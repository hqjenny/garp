module ConfigAddrDecoder(
    input [4:0] io_addr,
    output[31:0] io_en
);

  wire[31:0] T288;
  wire[32:0] T0;
  wire[32:0] T289;
  wire[31:0] T1;
  wire[31:0] T290;
  wire[30:0] T2;
  wire[30:0] T291;
  wire[29:0] T3;
  wire[29:0] T292;
  wire[28:0] T4;
  wire[28:0] T293;
  wire[27:0] T5;
  wire[27:0] T294;
  wire[26:0] T6;
  wire[26:0] T295;
  wire[25:0] T7;
  wire[25:0] T296;
  wire[24:0] T8;
  wire[24:0] T297;
  wire[23:0] T9;
  wire[23:0] T298;
  wire[22:0] T10;
  wire[22:0] T299;
  wire[21:0] T11;
  wire[21:0] T300;
  wire[20:0] T12;
  wire[20:0] T301;
  wire[19:0] T13;
  wire[19:0] T302;
  wire[18:0] T14;
  wire[18:0] T303;
  wire[17:0] T15;
  wire[17:0] T304;
  wire[16:0] T16;
  wire[16:0] T305;
  wire[15:0] T17;
  wire[15:0] T306;
  wire[14:0] T18;
  wire[14:0] T307;
  wire[13:0] T19;
  wire[13:0] T308;
  wire[12:0] T20;
  wire[12:0] T309;
  wire[11:0] T21;
  wire[11:0] T310;
  wire[10:0] T22;
  wire[10:0] T311;
  wire[9:0] T23;
  wire[9:0] T312;
  wire[8:0] T24;
  wire[8:0] T313;
  wire[7:0] T25;
  wire[7:0] T314;
  wire[6:0] T26;
  wire[6:0] T315;
  wire[5:0] T27;
  wire[5:0] T316;
  wire[4:0] T28;
  wire[4:0] T317;
  wire[3:0] T29;
  wire[3:0] T318;
  wire[2:0] T30;
  wire[2:0] T319;
  wire[1:0] T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T320;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire[2:0] T40;
  wire[2:0] T41;
  wire[2:0] T42;
  wire[2:0] T321;
  wire T43;
  wire T44;
  wire[2:0] T45;
  wire[2:0] T46;
  wire[2:0] T322;
  wire T47;
  wire[3:0] T48;
  wire[3:0] T49;
  wire[3:0] T50;
  wire[3:0] T323;
  wire T51;
  wire T52;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T324;
  wire T55;
  wire[4:0] T56;
  wire[4:0] T57;
  wire[4:0] T58;
  wire[4:0] T325;
  wire T59;
  wire T60;
  wire[4:0] T61;
  wire[4:0] T62;
  wire[4:0] T326;
  wire T63;
  wire[5:0] T64;
  wire[5:0] T65;
  wire[5:0] T66;
  wire[5:0] T327;
  wire T67;
  wire T68;
  wire[5:0] T69;
  wire[5:0] T70;
  wire[5:0] T328;
  wire T71;
  wire[6:0] T72;
  wire[6:0] T73;
  wire[6:0] T74;
  wire[6:0] T329;
  wire T75;
  wire T76;
  wire[6:0] T77;
  wire[6:0] T78;
  wire[6:0] T330;
  wire T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T331;
  wire T83;
  wire T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T332;
  wire T87;
  wire[8:0] T88;
  wire[8:0] T89;
  wire[8:0] T90;
  wire[8:0] T333;
  wire T91;
  wire T92;
  wire[8:0] T93;
  wire[8:0] T94;
  wire[8:0] T334;
  wire T95;
  wire[9:0] T96;
  wire[9:0] T97;
  wire[9:0] T98;
  wire[9:0] T335;
  wire T99;
  wire T100;
  wire[9:0] T101;
  wire[9:0] T102;
  wire[9:0] T336;
  wire T103;
  wire[10:0] T104;
  wire[10:0] T105;
  wire[10:0] T106;
  wire[10:0] T337;
  wire T107;
  wire T108;
  wire[10:0] T109;
  wire[10:0] T110;
  wire[10:0] T338;
  wire T111;
  wire[11:0] T112;
  wire[11:0] T113;
  wire[11:0] T114;
  wire[11:0] T339;
  wire T115;
  wire T116;
  wire[11:0] T117;
  wire[11:0] T118;
  wire[11:0] T340;
  wire T119;
  wire[12:0] T120;
  wire[12:0] T121;
  wire[12:0] T122;
  wire[12:0] T341;
  wire T123;
  wire T124;
  wire[12:0] T125;
  wire[12:0] T126;
  wire[12:0] T342;
  wire T127;
  wire[13:0] T128;
  wire[13:0] T129;
  wire[13:0] T130;
  wire[13:0] T343;
  wire T131;
  wire T132;
  wire[13:0] T133;
  wire[13:0] T134;
  wire[13:0] T344;
  wire T135;
  wire[14:0] T136;
  wire[14:0] T137;
  wire[14:0] T138;
  wire[14:0] T345;
  wire T139;
  wire T140;
  wire[14:0] T141;
  wire[14:0] T142;
  wire[14:0] T346;
  wire T143;
  wire[15:0] T144;
  wire[15:0] T145;
  wire[15:0] T146;
  wire[15:0] T347;
  wire T147;
  wire T148;
  wire[15:0] T149;
  wire[15:0] T150;
  wire[15:0] T348;
  wire T151;
  wire[16:0] T152;
  wire[16:0] T153;
  wire[16:0] T154;
  wire[16:0] T349;
  wire T155;
  wire T156;
  wire[16:0] T157;
  wire[16:0] T158;
  wire[16:0] T350;
  wire T159;
  wire[17:0] T160;
  wire[17:0] T161;
  wire[17:0] T162;
  wire[17:0] T351;
  wire T163;
  wire T164;
  wire[17:0] T165;
  wire[17:0] T166;
  wire[17:0] T352;
  wire T167;
  wire[18:0] T168;
  wire[18:0] T169;
  wire[18:0] T170;
  wire[18:0] T353;
  wire T171;
  wire T172;
  wire[18:0] T173;
  wire[18:0] T174;
  wire[18:0] T354;
  wire T175;
  wire[19:0] T176;
  wire[19:0] T177;
  wire[19:0] T178;
  wire[19:0] T355;
  wire T179;
  wire T180;
  wire[19:0] T181;
  wire[19:0] T182;
  wire[19:0] T356;
  wire T183;
  wire[20:0] T184;
  wire[20:0] T185;
  wire[20:0] T186;
  wire[20:0] T357;
  wire T187;
  wire T188;
  wire[20:0] T189;
  wire[20:0] T190;
  wire[20:0] T358;
  wire T191;
  wire[21:0] T192;
  wire[21:0] T193;
  wire[21:0] T194;
  wire[21:0] T359;
  wire T195;
  wire T196;
  wire[21:0] T197;
  wire[21:0] T198;
  wire[21:0] T360;
  wire T199;
  wire[22:0] T200;
  wire[22:0] T201;
  wire[22:0] T202;
  wire[22:0] T361;
  wire T203;
  wire T204;
  wire[22:0] T205;
  wire[22:0] T206;
  wire[22:0] T362;
  wire T207;
  wire[23:0] T208;
  wire[23:0] T209;
  wire[23:0] T210;
  wire[23:0] T363;
  wire T211;
  wire T212;
  wire[23:0] T213;
  wire[23:0] T214;
  wire[23:0] T364;
  wire T215;
  wire[24:0] T216;
  wire[24:0] T217;
  wire[24:0] T218;
  wire[24:0] T365;
  wire T219;
  wire T220;
  wire[24:0] T221;
  wire[24:0] T222;
  wire[24:0] T366;
  wire T223;
  wire[25:0] T224;
  wire[25:0] T225;
  wire[25:0] T226;
  wire[25:0] T367;
  wire T227;
  wire T228;
  wire[25:0] T229;
  wire[25:0] T230;
  wire[25:0] T368;
  wire T231;
  wire[26:0] T232;
  wire[26:0] T233;
  wire[26:0] T234;
  wire[26:0] T369;
  wire T235;
  wire T236;
  wire[26:0] T237;
  wire[26:0] T238;
  wire[26:0] T370;
  wire T239;
  wire[27:0] T240;
  wire[27:0] T241;
  wire[27:0] T242;
  wire[27:0] T371;
  wire T243;
  wire T244;
  wire[27:0] T245;
  wire[27:0] T246;
  wire[27:0] T372;
  wire T247;
  wire[28:0] T248;
  wire[28:0] T249;
  wire[28:0] T250;
  wire[28:0] T373;
  wire T251;
  wire T252;
  wire[28:0] T253;
  wire[28:0] T254;
  wire[28:0] T374;
  wire T255;
  wire[29:0] T256;
  wire[29:0] T257;
  wire[29:0] T258;
  wire[29:0] T375;
  wire T259;
  wire T260;
  wire[29:0] T261;
  wire[29:0] T262;
  wire[29:0] T376;
  wire T263;
  wire[30:0] T264;
  wire[30:0] T265;
  wire[30:0] T266;
  wire[30:0] T377;
  wire T267;
  wire T268;
  wire[30:0] T269;
  wire[30:0] T270;
  wire[30:0] T378;
  wire T271;
  wire[31:0] T272;
  wire[31:0] T273;
  wire[31:0] T274;
  wire[31:0] T379;
  wire T275;
  wire T276;
  wire[31:0] T277;
  wire[31:0] T278;
  wire[31:0] T380;
  wire T279;
  wire[32:0] T280;
  wire[32:0] T281;
  wire[32:0] T282;
  wire[32:0] T381;
  wire T283;
  wire T284;
  wire[32:0] T285;
  wire[32:0] T286;
  wire[32:0] T382;
  wire T287;


  assign io_en = T288;
  assign T288 = T0[5'h1f:1'h0];
  assign T0 = T287 ? T280 : T289;
  assign T289 = {1'h0, T1};
  assign T1 = T279 ? T272 : T290;
  assign T290 = {1'h0, T2};
  assign T2 = T271 ? T264 : T291;
  assign T291 = {1'h0, T3};
  assign T3 = T263 ? T256 : T292;
  assign T292 = {1'h0, T4};
  assign T4 = T255 ? T248 : T293;
  assign T293 = {1'h0, T5};
  assign T5 = T247 ? T240 : T294;
  assign T294 = {1'h0, T6};
  assign T6 = T239 ? T232 : T295;
  assign T295 = {1'h0, T7};
  assign T7 = T231 ? T224 : T296;
  assign T296 = {1'h0, T8};
  assign T8 = T223 ? T216 : T297;
  assign T297 = {1'h0, T9};
  assign T9 = T215 ? T208 : T298;
  assign T298 = {1'h0, T10};
  assign T10 = T207 ? T200 : T299;
  assign T299 = {1'h0, T11};
  assign T11 = T199 ? T192 : T300;
  assign T300 = {1'h0, T12};
  assign T12 = T191 ? T184 : T301;
  assign T301 = {1'h0, T13};
  assign T13 = T183 ? T176 : T302;
  assign T302 = {1'h0, T14};
  assign T14 = T175 ? T168 : T303;
  assign T303 = {1'h0, T15};
  assign T15 = T167 ? T160 : T304;
  assign T304 = {1'h0, T16};
  assign T16 = T159 ? T152 : T305;
  assign T305 = {1'h0, T17};
  assign T17 = T151 ? T144 : T306;
  assign T306 = {1'h0, T18};
  assign T18 = T143 ? T136 : T307;
  assign T307 = {1'h0, T19};
  assign T19 = T135 ? T128 : T308;
  assign T308 = {1'h0, T20};
  assign T20 = T127 ? T120 : T309;
  assign T309 = {1'h0, T21};
  assign T21 = T119 ? T112 : T310;
  assign T310 = {1'h0, T22};
  assign T22 = T111 ? T104 : T311;
  assign T311 = {1'h0, T23};
  assign T23 = T103 ? T96 : T312;
  assign T312 = {1'h0, T24};
  assign T24 = T95 ? T88 : T313;
  assign T313 = {1'h0, T25};
  assign T25 = T87 ? T80 : T314;
  assign T314 = {1'h0, T26};
  assign T26 = T79 ? T72 : T315;
  assign T315 = {1'h0, T27};
  assign T27 = T71 ? T64 : T316;
  assign T316 = {1'h0, T28};
  assign T28 = T63 ? T56 : T317;
  assign T317 = {1'h0, T29};
  assign T29 = T55 ? T48 : T318;
  assign T318 = {1'h0, T30};
  assign T30 = T47 ? T40 : T319;
  assign T319 = {1'h0, T31};
  assign T31 = T39 ? T32 : 2'h0;
  assign T32 = T37 | T33;
  assign T33 = T320 & T34;
  assign T34 = 2'h1;
  assign T320 = T35 ? 2'h3 : 2'h0;
  assign T35 = T36;
  assign T36 = 1'h1;
  assign T37 = 2'h0 & T38;
  assign T38 = ~ T34;
  assign T39 = io_addr == 5'h0;
  assign T40 = T45 | T41;
  assign T41 = T321 & T42;
  assign T42 = 3'h2;
  assign T321 = T43 ? 3'h7 : 3'h0;
  assign T43 = T44;
  assign T44 = 1'h1;
  assign T45 = T322 & T46;
  assign T46 = ~ T42;
  assign T322 = {1'h0, T31};
  assign T47 = io_addr == 5'h1;
  assign T48 = T53 | T49;
  assign T49 = T323 & T50;
  assign T50 = 4'h4;
  assign T323 = T51 ? 4'hf : 4'h0;
  assign T51 = T52;
  assign T52 = 1'h1;
  assign T53 = T324 & T54;
  assign T54 = ~ T50;
  assign T324 = {1'h0, T30};
  assign T55 = io_addr == 5'h2;
  assign T56 = T61 | T57;
  assign T57 = T325 & T58;
  assign T58 = 5'h8;
  assign T325 = T59 ? 5'h1f : 5'h0;
  assign T59 = T60;
  assign T60 = 1'h1;
  assign T61 = T326 & T62;
  assign T62 = ~ T58;
  assign T326 = {1'h0, T29};
  assign T63 = io_addr == 5'h3;
  assign T64 = T69 | T65;
  assign T65 = T327 & T66;
  assign T66 = 6'h10;
  assign T327 = T67 ? 6'h3f : 6'h0;
  assign T67 = T68;
  assign T68 = 1'h1;
  assign T69 = T328 & T70;
  assign T70 = ~ T66;
  assign T328 = {1'h0, T28};
  assign T71 = io_addr == 5'h4;
  assign T72 = T77 | T73;
  assign T73 = T329 & T74;
  assign T74 = 7'h20;
  assign T329 = T75 ? 7'h7f : 7'h0;
  assign T75 = T76;
  assign T76 = 1'h1;
  assign T77 = T330 & T78;
  assign T78 = ~ T74;
  assign T330 = {1'h0, T27};
  assign T79 = io_addr == 5'h5;
  assign T80 = T85 | T81;
  assign T81 = T331 & T82;
  assign T82 = 8'h40;
  assign T331 = T83 ? 8'hff : 8'h0;
  assign T83 = T84;
  assign T84 = 1'h1;
  assign T85 = T332 & T86;
  assign T86 = ~ T82;
  assign T332 = {1'h0, T26};
  assign T87 = io_addr == 5'h6;
  assign T88 = T93 | T89;
  assign T89 = T333 & T90;
  assign T90 = 9'h80;
  assign T333 = T91 ? 9'h1ff : 9'h0;
  assign T91 = T92;
  assign T92 = 1'h1;
  assign T93 = T334 & T94;
  assign T94 = ~ T90;
  assign T334 = {1'h0, T25};
  assign T95 = io_addr == 5'h7;
  assign T96 = T101 | T97;
  assign T97 = T335 & T98;
  assign T98 = 10'h100;
  assign T335 = T99 ? 10'h3ff : 10'h0;
  assign T99 = T100;
  assign T100 = 1'h1;
  assign T101 = T336 & T102;
  assign T102 = ~ T98;
  assign T336 = {1'h0, T24};
  assign T103 = io_addr == 5'h8;
  assign T104 = T109 | T105;
  assign T105 = T337 & T106;
  assign T106 = 11'h200;
  assign T337 = T107 ? 11'h7ff : 11'h0;
  assign T107 = T108;
  assign T108 = 1'h1;
  assign T109 = T338 & T110;
  assign T110 = ~ T106;
  assign T338 = {1'h0, T23};
  assign T111 = io_addr == 5'h9;
  assign T112 = T117 | T113;
  assign T113 = T339 & T114;
  assign T114 = 12'h400;
  assign T339 = T115 ? 12'hfff : 12'h0;
  assign T115 = T116;
  assign T116 = 1'h1;
  assign T117 = T340 & T118;
  assign T118 = ~ T114;
  assign T340 = {1'h0, T22};
  assign T119 = io_addr == 5'ha;
  assign T120 = T125 | T121;
  assign T121 = T341 & T122;
  assign T122 = 13'h800;
  assign T341 = T123 ? 13'h1fff : 13'h0;
  assign T123 = T124;
  assign T124 = 1'h1;
  assign T125 = T342 & T126;
  assign T126 = ~ T122;
  assign T342 = {1'h0, T21};
  assign T127 = io_addr == 5'hb;
  assign T128 = T133 | T129;
  assign T129 = T343 & T130;
  assign T130 = 14'h1000;
  assign T343 = T131 ? 14'h3fff : 14'h0;
  assign T131 = T132;
  assign T132 = 1'h1;
  assign T133 = T344 & T134;
  assign T134 = ~ T130;
  assign T344 = {1'h0, T20};
  assign T135 = io_addr == 5'hc;
  assign T136 = T141 | T137;
  assign T137 = T345 & T138;
  assign T138 = 15'h2000;
  assign T345 = T139 ? 15'h7fff : 15'h0;
  assign T139 = T140;
  assign T140 = 1'h1;
  assign T141 = T346 & T142;
  assign T142 = ~ T138;
  assign T346 = {1'h0, T19};
  assign T143 = io_addr == 5'hd;
  assign T144 = T149 | T145;
  assign T145 = T347 & T146;
  assign T146 = 16'h4000;
  assign T347 = T147 ? 16'hffff : 16'h0;
  assign T147 = T148;
  assign T148 = 1'h1;
  assign T149 = T348 & T150;
  assign T150 = ~ T146;
  assign T348 = {1'h0, T18};
  assign T151 = io_addr == 5'he;
  assign T152 = T157 | T153;
  assign T153 = T349 & T154;
  assign T154 = 17'h8000;
  assign T349 = T155 ? 17'h1ffff : 17'h0;
  assign T155 = T156;
  assign T156 = 1'h1;
  assign T157 = T350 & T158;
  assign T158 = ~ T154;
  assign T350 = {1'h0, T17};
  assign T159 = io_addr == 5'hf;
  assign T160 = T165 | T161;
  assign T161 = T351 & T162;
  assign T162 = 18'h10000;
  assign T351 = T163 ? 18'h3ffff : 18'h0;
  assign T163 = T164;
  assign T164 = 1'h1;
  assign T165 = T352 & T166;
  assign T166 = ~ T162;
  assign T352 = {1'h0, T16};
  assign T167 = io_addr == 5'h10;
  assign T168 = T173 | T169;
  assign T169 = T353 & T170;
  assign T170 = 19'h20000;
  assign T353 = T171 ? 19'h7ffff : 19'h0;
  assign T171 = T172;
  assign T172 = 1'h1;
  assign T173 = T354 & T174;
  assign T174 = ~ T170;
  assign T354 = {1'h0, T15};
  assign T175 = io_addr == 5'h11;
  assign T176 = T181 | T177;
  assign T177 = T355 & T178;
  assign T178 = 20'h40000;
  assign T355 = T179 ? 20'hfffff : 20'h0;
  assign T179 = T180;
  assign T180 = 1'h1;
  assign T181 = T356 & T182;
  assign T182 = ~ T178;
  assign T356 = {1'h0, T14};
  assign T183 = io_addr == 5'h12;
  assign T184 = T189 | T185;
  assign T185 = T357 & T186;
  assign T186 = 21'h80000;
  assign T357 = T187 ? 21'h1fffff : 21'h0;
  assign T187 = T188;
  assign T188 = 1'h1;
  assign T189 = T358 & T190;
  assign T190 = ~ T186;
  assign T358 = {1'h0, T13};
  assign T191 = io_addr == 5'h13;
  assign T192 = T197 | T193;
  assign T193 = T359 & T194;
  assign T194 = 22'h100000;
  assign T359 = T195 ? 22'h3fffff : 22'h0;
  assign T195 = T196;
  assign T196 = 1'h1;
  assign T197 = T360 & T198;
  assign T198 = ~ T194;
  assign T360 = {1'h0, T12};
  assign T199 = io_addr == 5'h14;
  assign T200 = T205 | T201;
  assign T201 = T361 & T202;
  assign T202 = 23'h200000;
  assign T361 = T203 ? 23'h7fffff : 23'h0;
  assign T203 = T204;
  assign T204 = 1'h1;
  assign T205 = T362 & T206;
  assign T206 = ~ T202;
  assign T362 = {1'h0, T11};
  assign T207 = io_addr == 5'h15;
  assign T208 = T213 | T209;
  assign T209 = T363 & T210;
  assign T210 = 24'h400000;
  assign T363 = T211 ? 24'hffffff : 24'h0;
  assign T211 = T212;
  assign T212 = 1'h1;
  assign T213 = T364 & T214;
  assign T214 = ~ T210;
  assign T364 = {1'h0, T10};
  assign T215 = io_addr == 5'h16;
  assign T216 = T221 | T217;
  assign T217 = T365 & T218;
  assign T218 = 25'h800000;
  assign T365 = T219 ? 25'h1ffffff : 25'h0;
  assign T219 = T220;
  assign T220 = 1'h1;
  assign T221 = T366 & T222;
  assign T222 = ~ T218;
  assign T366 = {1'h0, T9};
  assign T223 = io_addr == 5'h17;
  assign T224 = T229 | T225;
  assign T225 = T367 & T226;
  assign T226 = 26'h1000000;
  assign T367 = T227 ? 26'h3ffffff : 26'h0;
  assign T227 = T228;
  assign T228 = 1'h1;
  assign T229 = T368 & T230;
  assign T230 = ~ T226;
  assign T368 = {1'h0, T8};
  assign T231 = io_addr == 5'h18;
  assign T232 = T237 | T233;
  assign T233 = T369 & T234;
  assign T234 = 27'h2000000;
  assign T369 = T235 ? 27'h7ffffff : 27'h0;
  assign T235 = T236;
  assign T236 = 1'h1;
  assign T237 = T370 & T238;
  assign T238 = ~ T234;
  assign T370 = {1'h0, T7};
  assign T239 = io_addr == 5'h19;
  assign T240 = T245 | T241;
  assign T241 = T371 & T242;
  assign T242 = 28'h4000000;
  assign T371 = T243 ? 28'hfffffff : 28'h0;
  assign T243 = T244;
  assign T244 = 1'h1;
  assign T245 = T372 & T246;
  assign T246 = ~ T242;
  assign T372 = {1'h0, T6};
  assign T247 = io_addr == 5'h1a;
  assign T248 = T253 | T249;
  assign T249 = T373 & T250;
  assign T250 = 29'h8000000;
  assign T373 = T251 ? 29'h1fffffff : 29'h0;
  assign T251 = T252;
  assign T252 = 1'h1;
  assign T253 = T374 & T254;
  assign T254 = ~ T250;
  assign T374 = {1'h0, T5};
  assign T255 = io_addr == 5'h1b;
  assign T256 = T261 | T257;
  assign T257 = T375 & T258;
  assign T258 = 30'h10000000;
  assign T375 = T259 ? 30'h3fffffff : 30'h0;
  assign T259 = T260;
  assign T260 = 1'h1;
  assign T261 = T376 & T262;
  assign T262 = ~ T258;
  assign T376 = {1'h0, T4};
  assign T263 = io_addr == 5'h1c;
  assign T264 = T269 | T265;
  assign T265 = T377 & T266;
  assign T266 = 31'h20000000;
  assign T377 = T267 ? 31'h7fffffff : 31'h0;
  assign T267 = T268;
  assign T268 = 1'h1;
  assign T269 = T378 & T270;
  assign T270 = ~ T266;
  assign T378 = {1'h0, T3};
  assign T271 = io_addr == 5'h1d;
  assign T272 = T277 | T273;
  assign T273 = T379 & T274;
  assign T274 = 32'h40000000;
  assign T379 = T275 ? 32'hffffffff : 32'h0;
  assign T275 = T276;
  assign T276 = 1'h1;
  assign T277 = T380 & T278;
  assign T278 = ~ T274;
  assign T380 = {1'h0, T2};
  assign T279 = io_addr == 5'h1e;
  assign T280 = T285 | T281;
  assign T281 = T381 & T282;
  assign T282 = 33'h80000000;
  assign T381 = T283 ? 33'h1ffffffff : 33'h0;
  assign T283 = T284;
  assign T284 = 1'h1;
  assign T285 = T382 & T286;
  assign T286 = ~ T282;
  assign T382 = {1'h0, T1};
  assign T287 = io_addr == 5'h1f;
endmodule

module ConfigurationModule(input clk, input reset,
    input [1:0] io_in,
    input  io_en,
    output[63:0] io_out
);

  reg [63:0] config_reg;
  wire[63:0] T21;
  wire[64:0] T22;
  wire[64:0] T0;
  wire[64:0] T1;
  wire[64:0] T23;
  wire[63:0] T2;
  wire[63:0] T24;
  wire[61:0] T3;
  wire[64:0] T4;
  wire[64:0] T5;
  wire[64:0] T6;
  wire[64:0] T25;
  wire T7;
  wire T8;
  wire T9;
  wire[64:0] T10;
  wire[64:0] T11;
  wire[64:0] T26;
  wire[64:0] T12;
  wire[64:0] T27;
  wire[63:0] T13;
  wire[63:0] T14;
  wire[63:0] T28;
  wire T15;
  wire T16;
  wire T17;
  wire T29;
  wire[64:0] T18;
  wire[64:0] T30;
  wire[63:0] T19;
  wire T31;
  wire T20;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    config_reg = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_out = config_reg;
  assign T21 = T22[6'h3f:1'h0];
  assign T22 = reset ? 65'h0 : T0;
  assign T0 = T20 ? T12 : T1;
  assign T1 = T20 ? T4 : T23;
  assign T23 = {1'h0, T2};
  assign T2 = T20 ? T24 : config_reg;
  assign T24 = {2'h0, T3};
  assign T3 = config_reg >> 2'h2;
  assign T4 = T10 | T5;
  assign T5 = T25 & T6;
  assign T6 = 65'h8000000000000000;
  assign T25 = T7 ? 65'h1ffffffffffffffff : 65'h0;
  assign T7 = T8;
  assign T8 = T9;
  assign T9 = io_in[1'h1];
  assign T10 = T26 & T11;
  assign T11 = ~ T6;
  assign T26 = {1'h0, T2};
  assign T12 = T18 | T27;
  assign T27 = {T29, T13};
  assign T13 = T28 & T14;
  assign T14 = 64'h4000000000000000;
  assign T28 = T15 ? 64'hffffffffffffffff : 64'h0;
  assign T15 = T16;
  assign T16 = T17;
  assign T17 = io_in[1'h0];
  assign T29 = T13[6'h3f];
  assign T18 = T1 & T30;
  assign T30 = {T31, T19};
  assign T19 = ~ T14;
  assign T31 = T19[6'h3f];
  assign T20 = io_en;

  always @(posedge clk) begin
    config_reg <= T21;
  end
endmodule

module ControlMuxModule(
    input [1:0] io_h_wire_above_8,
    input [1:0] io_h_wire_above_7,
    input [1:0] io_h_wire_above_6,
    input [1:0] io_h_wire_above_5,
    input [1:0] io_h_wire_above_4,
    input [1:0] io_h_wire_above_3,
    input [1:0] io_h_wire_above_2,
    input [1:0] io_h_wire_above_1,
    input [1:0] io_h_wire_above_0,
    input [1:0] io_h_wire_below_8,
    input [1:0] io_h_wire_below_7,
    input [1:0] io_h_wire_below_6,
    input [1:0] io_h_wire_below_5,
    input [1:0] io_h_wire_below_4,
    input [1:0] io_h_wire_below_3,
    input [1:0] io_h_wire_below_2,
    input [1:0] io_h_wire_below_1,
    input [1:0] io_h_wire_below_0,
    input [5:0] io_select,
    output[1:0] io_a
);

  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire[3:0] T18;
  wire T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[1:0] T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire[1:0] T35;
  wire T36;
  wire T37;
  wire[1:0] T38;
  wire T39;
  wire T40;
  wire[1:0] T41;
  wire T42;
  wire T43;


  assign io_a = T0;
  assign T0 = T42 ? T41 : T1;
  assign T1 = T39 ? T38 : T2;
  assign T2 = T36 ? T35 : T3;
  assign T3 = T33 ? T32 : T4;
  assign T4 = T30 ? T29 : T5;
  assign T5 = T27 ? T26 : T6;
  assign T6 = T24 ? T23 : T7;
  assign T7 = T21 ? T20 : T8;
  assign T8 = T16 ? T14 : T9;
  assign T9 = T12 ? T10 : 2'h0;
  assign T10 = {T11, 1'h0};
  assign T11 = io_select[1'h0];
  assign T12 = T13 == 1'h0;
  assign T13 = io_select[3'h5];
  assign T14 = T15 ? io_h_wire_below_0 : io_h_wire_above_0;
  assign T15 = io_select[3'h4];
  assign T16 = T19 & T17;
  assign T17 = 4'h2 == T18;
  assign T18 = io_select[2'h3:1'h0];
  assign T19 = T12 ^ 1'h1;
  assign T20 = T15 ? io_h_wire_below_1 : io_h_wire_above_1;
  assign T21 = T19 & T22;
  assign T22 = 4'h3 == T18;
  assign T23 = T15 ? io_h_wire_below_2 : io_h_wire_above_2;
  assign T24 = T19 & T25;
  assign T25 = 4'h4 == T18;
  assign T26 = T15 ? io_h_wire_below_3 : io_h_wire_above_3;
  assign T27 = T19 & T28;
  assign T28 = 4'h5 == T18;
  assign T29 = T15 ? io_h_wire_below_4 : io_h_wire_above_4;
  assign T30 = T19 & T31;
  assign T31 = 4'h6 == T18;
  assign T32 = T15 ? io_h_wire_below_5 : io_h_wire_above_5;
  assign T33 = T19 & T34;
  assign T34 = 4'h7 == T18;
  assign T35 = T15 ? io_h_wire_below_6 : io_h_wire_above_6;
  assign T36 = T19 & T37;
  assign T37 = 4'h8 == T18;
  assign T38 = T15 ? io_h_wire_below_7 : io_h_wire_above_7;
  assign T39 = T19 & T40;
  assign T40 = 4'h9 == T18;
  assign T41 = T15 ? io_h_wire_below_8 : io_h_wire_above_8;
  assign T42 = T19 & T43;
  assign T43 = 4'ha == T18;
endmodule

module ControlReducerModule(
    input [1:0] io_a,
    input [1:0] io_select,
    output io_out
);

  wire T0;
  wire T1;
  wire T2;
  wire a0;
  wire T3;
  wire a1;
  wire T4;
  wire T5;
  wire T6;


  assign io_out = T0;
  assign T0 = T4 ? a1 : T1;
  assign T1 = T3 ? a0 : T2;
  assign T2 = a0 | a1;
  assign a0 = io_a[1'h0];
  assign T3 = io_select == 2'h0;
  assign a1 = io_a[1'h1];
  assign T4 = T6 & T5;
  assign T5 = io_select == 2'h3;
  assign T6 = T3 ^ 1'h1;
endmodule

module ControlBlockModule(input clk, input reset,
    input [1:0] io_H_wire_above_in_8,
    input [1:0] io_H_wire_above_in_7,
    input [1:0] io_H_wire_above_in_6,
    input [1:0] io_H_wire_above_in_5,
    input [1:0] io_H_wire_above_in_4,
    input [1:0] io_H_wire_above_in_3,
    input [1:0] io_H_wire_above_in_2,
    input [1:0] io_H_wire_above_in_1,
    input [1:0] io_H_wire_above_in_0,
    input [1:0] io_H_wire_below_in_8,
    input [1:0] io_H_wire_below_in_7,
    input [1:0] io_H_wire_below_in_6,
    input [1:0] io_H_wire_below_in_5,
    input [1:0] io_H_wire_below_in_4,
    input [1:0] io_H_wire_below_in_3,
    input [1:0] io_H_wire_below_in_2,
    input [1:0] io_H_wire_below_in_1,
    input [1:0] io_H_wire_below_in_0,
    input [63:0] io_config,
    output[1:0] io_Hdir,
    output io_read_demand_access,
    output io_write_demand_access,
    output io_prefetch_demand_access,
    output io_load_transfer_access,
    output io_store_transfer_access,
    output io_mem_D_or_Z
);

  reg  T0;
  wire T1;
  wire T2;
  wire[1:0] bus;
  wire[1:0] T3;
  reg  T4;
  wire T5;
  wire T6;
  wire[1:0] K;
  wire[1:0] T7;
  wire[1:0] primes_3;
  wire[1:0] T8;
  wire[1:0] primes_2;
  wire[1:0] T9;
  wire[1:0] primes_1;
  wire[1:0] T10;
  wire[1:0] primes_0;
  wire[1:0] T11;
  wire[5:0] indexes_3;
  wire[5:0] T12;
  wire[5:0] indexes_2;
  wire[5:0] T13;
  wire[5:0] indexes_1;
  wire[5:0] T14;
  wire[5:0] indexes_0;
  wire[5:0] T15;
  wire R;
  wire T16;
  wire T17;
  wire D_prime;
  wire T18;
  wire T19;
  wire transfer_access;
  wire T20;
  wire C_prime;
  wire T21;
  wire T22;
  wire T23;
  wire A_prime;
  wire T24;
  wire mem_mode;
  wire T25;
  wire[2:0] mode;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[1:0] demand_access_type;
  wire[1:0] T32;
  wire T33;
  wire demand_access;
  wire T34;
  wire B_prime;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] ControlMuxModule_io_a;
  wire[1:0] ControlMuxModule_1_io_a;
  wire[1:0] ControlMuxModule_2_io_a;
  wire[1:0] ControlMuxModule_3_io_a;
  wire ControlReducerModule_io_out;
  wire ControlReducerModule_1_io_out;
  wire ControlReducerModule_2_io_out;
  wire ControlReducerModule_3_io_out;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    T4 = 1'b0;
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = bus == 2'h0;
  assign bus = T3;
  assign T3 = io_config[4'h9:4'h8];
  assign T5 = T6 | reset;
  assign T6 = K == 2'h0;
  assign K = T7;
  assign T7 = io_config[5'h11:5'h10];
  assign primes_3 = T8;
  assign T8 = io_config[6'h21:6'h20];
  assign primes_2 = T9;
  assign T9 = io_config[6'h29:6'h28];
  assign primes_1 = T10;
  assign T10 = io_config[6'h31:6'h30];
  assign primes_0 = T11;
  assign T11 = io_config[6'h39:6'h38];
  assign indexes_3 = T12;
  assign T12 = io_config[6'h27:6'h22];
  assign indexes_2 = T13;
  assign T13 = io_config[6'h2f:6'h2a];
  assign indexes_1 = T14;
  assign T14 = io_config[6'h37:6'h32];
  assign indexes_0 = T15;
  assign T15 = io_config[6'h3f:6'h3a];
  assign io_mem_D_or_Z = R;
  assign R = T16;
  assign T16 = io_config[4'hd];
  assign io_store_transfer_access = T17;
  assign T17 = transfer_access & D_prime;
  assign D_prime = T18;
  assign T18 = T19;
  assign T19 = ControlReducerModule_io_out & ControlReducerModule_3_io_out;
  assign transfer_access = T20;
  assign T20 = T23 & C_prime;
  assign C_prime = T21;
  assign T21 = T22;
  assign T22 = ControlReducerModule_io_out & ControlReducerModule_2_io_out;
  assign T23 = mem_mode & A_prime;
  assign A_prime = T24;
  assign T24 = ControlReducerModule_io_out;
  assign mem_mode = T25;
  assign T25 = mode == 3'h6;
  assign mode = io_config[2'h2:1'h0];
  assign io_load_transfer_access = T26;
  assign T26 = transfer_access & T27;
  assign T27 = ~ D_prime;
  assign io_prefetch_demand_access = T28;
  assign T28 = T33 & T29;
  assign T29 = ~ T30;
  assign T30 = T31;
  assign T31 = demand_access_type[1'h1];
  assign demand_access_type = T32;
  assign T32 = io_config[5'h1f:5'h1e];
  assign T33 = demand_access & D_prime;
  assign demand_access = T34;
  assign T34 = T37 & B_prime;
  assign B_prime = T35;
  assign T35 = T36;
  assign T36 = ControlReducerModule_io_out & ControlReducerModule_1_io_out;
  assign T37 = mem_mode & A_prime;
  assign io_write_demand_access = T38;
  assign T38 = T41 & T39;
  assign T39 = T40;
  assign T40 = demand_access_type[1'h1];
  assign T41 = demand_access & D_prime;
  assign io_read_demand_access = T42;
  assign T42 = demand_access & T43;
  assign T43 = ~ D_prime;
  assign io_Hdir = T44;
  assign T44 = io_config[3'h4:2'h3];
  ControlMuxModule ControlMuxModule(
       .io_h_wire_above_8( io_H_wire_above_in_8 ),
       .io_h_wire_above_7( io_H_wire_above_in_7 ),
       .io_h_wire_above_6( io_H_wire_above_in_6 ),
       .io_h_wire_above_5( io_H_wire_above_in_5 ),
       .io_h_wire_above_4( io_H_wire_above_in_4 ),
       .io_h_wire_above_3( io_H_wire_above_in_3 ),
       .io_h_wire_above_2( io_H_wire_above_in_2 ),
       .io_h_wire_above_1( io_H_wire_above_in_1 ),
       .io_h_wire_above_0( io_H_wire_above_in_0 ),
       .io_h_wire_below_8( io_H_wire_below_in_8 ),
       .io_h_wire_below_7( io_H_wire_below_in_7 ),
       .io_h_wire_below_6( io_H_wire_below_in_6 ),
       .io_h_wire_below_5( io_H_wire_below_in_5 ),
       .io_h_wire_below_4( io_H_wire_below_in_4 ),
       .io_h_wire_below_3( io_H_wire_below_in_3 ),
       .io_h_wire_below_2( io_H_wire_below_in_2 ),
       .io_h_wire_below_1( io_H_wire_below_in_1 ),
       .io_h_wire_below_0( io_H_wire_below_in_0 ),
       .io_select( indexes_0 ),
       .io_a( ControlMuxModule_io_a )
  );
  ControlMuxModule ControlMuxModule_1(
       .io_h_wire_above_8( io_H_wire_above_in_8 ),
       .io_h_wire_above_7( io_H_wire_above_in_7 ),
       .io_h_wire_above_6( io_H_wire_above_in_6 ),
       .io_h_wire_above_5( io_H_wire_above_in_5 ),
       .io_h_wire_above_4( io_H_wire_above_in_4 ),
       .io_h_wire_above_3( io_H_wire_above_in_3 ),
       .io_h_wire_above_2( io_H_wire_above_in_2 ),
       .io_h_wire_above_1( io_H_wire_above_in_1 ),
       .io_h_wire_above_0( io_H_wire_above_in_0 ),
       .io_h_wire_below_8( io_H_wire_below_in_8 ),
       .io_h_wire_below_7( io_H_wire_below_in_7 ),
       .io_h_wire_below_6( io_H_wire_below_in_6 ),
       .io_h_wire_below_5( io_H_wire_below_in_5 ),
       .io_h_wire_below_4( io_H_wire_below_in_4 ),
       .io_h_wire_below_3( io_H_wire_below_in_3 ),
       .io_h_wire_below_2( io_H_wire_below_in_2 ),
       .io_h_wire_below_1( io_H_wire_below_in_1 ),
       .io_h_wire_below_0( io_H_wire_below_in_0 ),
       .io_select( indexes_1 ),
       .io_a( ControlMuxModule_1_io_a )
  );
  ControlMuxModule ControlMuxModule_2(
       .io_h_wire_above_8( io_H_wire_above_in_8 ),
       .io_h_wire_above_7( io_H_wire_above_in_7 ),
       .io_h_wire_above_6( io_H_wire_above_in_6 ),
       .io_h_wire_above_5( io_H_wire_above_in_5 ),
       .io_h_wire_above_4( io_H_wire_above_in_4 ),
       .io_h_wire_above_3( io_H_wire_above_in_3 ),
       .io_h_wire_above_2( io_H_wire_above_in_2 ),
       .io_h_wire_above_1( io_H_wire_above_in_1 ),
       .io_h_wire_above_0( io_H_wire_above_in_0 ),
       .io_h_wire_below_8( io_H_wire_below_in_8 ),
       .io_h_wire_below_7( io_H_wire_below_in_7 ),
       .io_h_wire_below_6( io_H_wire_below_in_6 ),
       .io_h_wire_below_5( io_H_wire_below_in_5 ),
       .io_h_wire_below_4( io_H_wire_below_in_4 ),
       .io_h_wire_below_3( io_H_wire_below_in_3 ),
       .io_h_wire_below_2( io_H_wire_below_in_2 ),
       .io_h_wire_below_1( io_H_wire_below_in_1 ),
       .io_h_wire_below_0( io_H_wire_below_in_0 ),
       .io_select( indexes_2 ),
       .io_a( ControlMuxModule_2_io_a )
  );
  ControlMuxModule ControlMuxModule_3(
       .io_h_wire_above_8( io_H_wire_above_in_8 ),
       .io_h_wire_above_7( io_H_wire_above_in_7 ),
       .io_h_wire_above_6( io_H_wire_above_in_6 ),
       .io_h_wire_above_5( io_H_wire_above_in_5 ),
       .io_h_wire_above_4( io_H_wire_above_in_4 ),
       .io_h_wire_above_3( io_H_wire_above_in_3 ),
       .io_h_wire_above_2( io_H_wire_above_in_2 ),
       .io_h_wire_above_1( io_H_wire_above_in_1 ),
       .io_h_wire_above_0( io_H_wire_above_in_0 ),
       .io_h_wire_below_8( io_H_wire_below_in_8 ),
       .io_h_wire_below_7( io_H_wire_below_in_7 ),
       .io_h_wire_below_6( io_H_wire_below_in_6 ),
       .io_h_wire_below_5( io_H_wire_below_in_5 ),
       .io_h_wire_below_4( io_H_wire_below_in_4 ),
       .io_h_wire_below_3( io_H_wire_below_in_3 ),
       .io_h_wire_below_2( io_H_wire_below_in_2 ),
       .io_h_wire_below_1( io_H_wire_below_in_1 ),
       .io_h_wire_below_0( io_H_wire_below_in_0 ),
       .io_select( indexes_3 ),
       .io_a( ControlMuxModule_3_io_a )
  );
  ControlReducerModule ControlReducerModule(
       .io_a( ControlMuxModule_io_a ),
       .io_select( primes_0 ),
       .io_out( ControlReducerModule_io_out )
  );
  ControlReducerModule ControlReducerModule_1(
       .io_a( ControlMuxModule_1_io_a ),
       .io_select( primes_1 ),
       .io_out( ControlReducerModule_1_io_out )
  );
  ControlReducerModule ControlReducerModule_2(
       .io_a( ControlMuxModule_2_io_a ),
       .io_select( primes_2 ),
       .io_out( ControlReducerModule_2_io_out )
  );
  ControlReducerModule ControlReducerModule_3(
       .io_a( ControlMuxModule_3_io_a ),
       .io_select( primes_3 ),
       .io_out( ControlReducerModule_3_io_out )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T4 <= 1'b1;
  if(!T5 && T4 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "We only have 1 memory bus!\n");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "We only have memory bus 0!\n");
    $finish;
  end
// synthesis translate_on
`endif
  end
endmodule

module LogicBlockInBBModule(
    input [1:0] io_V_wire_in_15,
    input [1:0] io_V_wire_in_14,
    input [1:0] io_V_wire_in_13,
    input [1:0] io_V_wire_in_12,
    input [1:0] io_V_wire_in_11,
    input [1:0] io_V_wire_in_10,
    input [1:0] io_V_wire_in_9,
    input [1:0] io_V_wire_in_8,
    input [1:0] io_V_wire_in_7,
    input [1:0] io_V_wire_in_6,
    input [1:0] io_V_wire_in_5,
    input [1:0] io_V_wire_in_4,
    input [1:0] io_V_wire_in_3,
    input [1:0] io_V_wire_in_2,
    input [1:0] io_V_wire_in_1,
    input [1:0] io_V_wire_in_0,
    input [1:0] io_H_wire_above_in_10,
    input [1:0] io_H_wire_above_in_9,
    input [1:0] io_H_wire_above_in_8,
    input [1:0] io_H_wire_above_in_7,
    input [1:0] io_H_wire_above_in_6,
    input [1:0] io_H_wire_above_in_5,
    input [1:0] io_H_wire_above_in_4,
    input [1:0] io_H_wire_above_in_3,
    input [1:0] io_H_wire_above_in_2,
    input [1:0] io_H_wire_above_in_1,
    input [1:0] io_H_wire_above_in_0,
    input [1:0] io_H_wire_below_in_10,
    input [1:0] io_H_wire_below_in_9,
    input [1:0] io_H_wire_below_in_8,
    input [1:0] io_H_wire_below_in_7,
    input [1:0] io_H_wire_below_in_6,
    input [1:0] io_H_wire_below_in_5,
    input [1:0] io_H_wire_below_in_4,
    input [1:0] io_H_wire_below_in_3,
    input [1:0] io_H_wire_below_in_2,
    input [1:0] io_H_wire_below_in_1,
    input [1:0] io_H_wire_below_in_0,
    input [1:0] io_G_wire_above_in_3,
    input [1:0] io_G_wire_above_in_2,
    input [1:0] io_G_wire_above_in_1,
    input [1:0] io_G_wire_above_in_0,
    input [1:0] io_G_wire_below_in_3,
    input [1:0] io_G_wire_below_in_2,
    input [1:0] io_G_wire_below_in_1,
    input [1:0] io_G_wire_below_in_0,
    input [5:0] io_config_X_in_3,
    input [5:0] io_config_X_in_2,
    input [5:0] io_config_X_in_1,
    input [5:0] io_config_X_in_0,
    input [1:0] io_Z_reg,
    input [1:0] io_D_reg,
    output[1:0] io_X_in_3,
    output[1:0] io_X_in_2,
    output[1:0] io_X_in_1,
    output[1:0] io_X_in_0
);

  wire[23:0] T304;
  wire[24:0] T0;
  wire[24:0] T305;
  wire[23:0] T1;
  wire[5:0] T2;
  wire[24:0] T3;
  wire[24:0] T4;
  wire[24:0] T5;
  wire[24:0] T306;
  wire[18:0] T6;
  wire[18:0] T307;
  wire[17:0] T7;
  wire[5:0] T8;
  wire[18:0] T9;
  wire[18:0] T10;
  wire[18:0] T11;
  wire[18:0] T308;
  wire[12:0] T12;
  wire[12:0] T309;
  wire[11:0] T13;
  wire[5:0] T14;
  wire[12:0] T15;
  wire[12:0] T16;
  wire[12:0] T17;
  wire[12:0] T310;
  wire[6:0] T18;
  wire[6:0] T311;
  wire[5:0] T19;
  wire[5:0] T20;
  wire[6:0] T21;
  wire[6:0] T22;
  wire[6:0] T23;
  wire[7:0] T312;
  wire[8:0] T24;
  wire[8:0] T313;
  wire[7:0] T25;
  wire[1:0] T26;
  wire[8:0] T27;
  wire[8:0] T28;
  wire[8:0] T29;
  wire[8:0] T314;
  wire[6:0] T30;
  wire[6:0] T315;
  wire[5:0] T31;
  wire[1:0] T32;
  wire[6:0] T33;
  wire[6:0] T34;
  wire[6:0] T35;
  wire[6:0] T316;
  wire[4:0] T36;
  wire[4:0] T317;
  wire[3:0] T37;
  wire[1:0] T38;
  wire[4:0] T39;
  wire[4:0] T40;
  wire[4:0] T41;
  wire[4:0] T318;
  wire[2:0] T42;
  wire[2:0] T319;
  wire[1:0] T43;
  wire[1:0] T44;
  wire[2:0] T45;
  wire[2:0] T46;
  wire[2:0] T47;
  wire[7:0] T320;
  wire[8:0] T48;
  wire[8:0] T321;
  wire[7:0] T49;
  wire[1:0] T50;
  wire[8:0] T51;
  wire[8:0] T52;
  wire[8:0] T53;
  wire[8:0] T322;
  wire[6:0] T54;
  wire[6:0] T323;
  wire[5:0] T55;
  wire[1:0] T56;
  wire[6:0] T57;
  wire[6:0] T58;
  wire[6:0] T59;
  wire[6:0] T324;
  wire[4:0] T60;
  wire[4:0] T325;
  wire[3:0] T61;
  wire[1:0] T62;
  wire[4:0] T63;
  wire[4:0] T64;
  wire[4:0] T65;
  wire[4:0] T326;
  wire[2:0] T66;
  wire[2:0] T327;
  wire[1:0] T67;
  wire[1:0] T68;
  wire[2:0] T69;
  wire[2:0] T70;
  wire[2:0] T71;
  wire[21:0] T328;
  wire[22:0] T72;
  wire[22:0] T329;
  wire[21:0] T73;
  wire[1:0] T74;
  wire[22:0] T75;
  wire[22:0] T76;
  wire[22:0] T77;
  wire[22:0] T330;
  wire[20:0] T78;
  wire[20:0] T331;
  wire[19:0] T79;
  wire[1:0] T80;
  wire[20:0] T81;
  wire[20:0] T82;
  wire[20:0] T83;
  wire[20:0] T332;
  wire[18:0] T84;
  wire[18:0] T333;
  wire[17:0] T85;
  wire[1:0] T86;
  wire[18:0] T87;
  wire[18:0] T88;
  wire[18:0] T89;
  wire[18:0] T334;
  wire[16:0] T90;
  wire[16:0] T335;
  wire[15:0] T91;
  wire[1:0] T92;
  wire[16:0] T93;
  wire[16:0] T94;
  wire[16:0] T95;
  wire[16:0] T336;
  wire[14:0] T96;
  wire[14:0] T337;
  wire[13:0] T97;
  wire[1:0] T98;
  wire[14:0] T99;
  wire[14:0] T100;
  wire[14:0] T101;
  wire[14:0] T338;
  wire[12:0] T102;
  wire[12:0] T339;
  wire[11:0] T103;
  wire[1:0] T104;
  wire[12:0] T105;
  wire[12:0] T106;
  wire[12:0] T107;
  wire[12:0] T340;
  wire[10:0] T108;
  wire[10:0] T341;
  wire[9:0] T109;
  wire[1:0] T110;
  wire[10:0] T111;
  wire[10:0] T112;
  wire[10:0] T113;
  wire[10:0] T342;
  wire[8:0] T114;
  wire[8:0] T343;
  wire[7:0] T115;
  wire[1:0] T116;
  wire[8:0] T117;
  wire[8:0] T118;
  wire[8:0] T119;
  wire[8:0] T344;
  wire[6:0] T120;
  wire[6:0] T345;
  wire[5:0] T121;
  wire[1:0] T122;
  wire[6:0] T123;
  wire[6:0] T124;
  wire[6:0] T125;
  wire[6:0] T346;
  wire[4:0] T126;
  wire[4:0] T347;
  wire[3:0] T127;
  wire[1:0] T128;
  wire[4:0] T129;
  wire[4:0] T130;
  wire[4:0] T131;
  wire[4:0] T348;
  wire[2:0] T132;
  wire[2:0] T349;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[2:0] T135;
  wire[2:0] T136;
  wire[2:0] T137;
  wire[21:0] T350;
  wire[22:0] T138;
  wire[22:0] T351;
  wire[21:0] T139;
  wire[1:0] T140;
  wire[22:0] T141;
  wire[22:0] T142;
  wire[22:0] T143;
  wire[22:0] T352;
  wire[20:0] T144;
  wire[20:0] T353;
  wire[19:0] T145;
  wire[1:0] T146;
  wire[20:0] T147;
  wire[20:0] T148;
  wire[20:0] T149;
  wire[20:0] T354;
  wire[18:0] T150;
  wire[18:0] T355;
  wire[17:0] T151;
  wire[1:0] T152;
  wire[18:0] T153;
  wire[18:0] T154;
  wire[18:0] T155;
  wire[18:0] T356;
  wire[16:0] T156;
  wire[16:0] T357;
  wire[15:0] T157;
  wire[1:0] T158;
  wire[16:0] T159;
  wire[16:0] T160;
  wire[16:0] T161;
  wire[16:0] T358;
  wire[14:0] T162;
  wire[14:0] T359;
  wire[13:0] T163;
  wire[1:0] T164;
  wire[14:0] T165;
  wire[14:0] T166;
  wire[14:0] T167;
  wire[14:0] T360;
  wire[12:0] T168;
  wire[12:0] T361;
  wire[11:0] T169;
  wire[1:0] T170;
  wire[12:0] T171;
  wire[12:0] T172;
  wire[12:0] T173;
  wire[12:0] T362;
  wire[10:0] T174;
  wire[10:0] T363;
  wire[9:0] T175;
  wire[1:0] T176;
  wire[10:0] T177;
  wire[10:0] T178;
  wire[10:0] T179;
  wire[10:0] T364;
  wire[8:0] T180;
  wire[8:0] T365;
  wire[7:0] T181;
  wire[1:0] T182;
  wire[8:0] T183;
  wire[8:0] T184;
  wire[8:0] T185;
  wire[8:0] T366;
  wire[6:0] T186;
  wire[6:0] T367;
  wire[5:0] T187;
  wire[1:0] T188;
  wire[6:0] T189;
  wire[6:0] T190;
  wire[6:0] T191;
  wire[6:0] T368;
  wire[4:0] T192;
  wire[4:0] T369;
  wire[3:0] T193;
  wire[1:0] T194;
  wire[4:0] T195;
  wire[4:0] T196;
  wire[4:0] T197;
  wire[4:0] T370;
  wire[2:0] T198;
  wire[2:0] T371;
  wire[1:0] T199;
  wire[1:0] T200;
  wire[2:0] T201;
  wire[2:0] T202;
  wire[2:0] T203;
  wire[31:0] T372;
  wire[32:0] T204;
  wire[32:0] T373;
  wire[31:0] T205;
  wire[1:0] T206;
  wire[32:0] T207;
  wire[32:0] T208;
  wire[32:0] T209;
  wire[32:0] T374;
  wire[30:0] T210;
  wire[30:0] T375;
  wire[29:0] T211;
  wire[1:0] T212;
  wire[30:0] T213;
  wire[30:0] T214;
  wire[30:0] T215;
  wire[30:0] T376;
  wire[28:0] T216;
  wire[28:0] T377;
  wire[27:0] T217;
  wire[1:0] T218;
  wire[28:0] T219;
  wire[28:0] T220;
  wire[28:0] T221;
  wire[28:0] T378;
  wire[26:0] T222;
  wire[26:0] T379;
  wire[25:0] T223;
  wire[1:0] T224;
  wire[26:0] T225;
  wire[26:0] T226;
  wire[26:0] T227;
  wire[26:0] T380;
  wire[24:0] T228;
  wire[24:0] T381;
  wire[23:0] T229;
  wire[1:0] T230;
  wire[24:0] T231;
  wire[24:0] T232;
  wire[24:0] T233;
  wire[24:0] T382;
  wire[22:0] T234;
  wire[22:0] T383;
  wire[21:0] T235;
  wire[1:0] T236;
  wire[22:0] T237;
  wire[22:0] T238;
  wire[22:0] T239;
  wire[22:0] T384;
  wire[20:0] T240;
  wire[20:0] T385;
  wire[19:0] T241;
  wire[1:0] T242;
  wire[20:0] T243;
  wire[20:0] T244;
  wire[20:0] T245;
  wire[20:0] T386;
  wire[18:0] T246;
  wire[18:0] T387;
  wire[17:0] T247;
  wire[1:0] T248;
  wire[18:0] T249;
  wire[18:0] T250;
  wire[18:0] T251;
  wire[18:0] T388;
  wire[16:0] T252;
  wire[16:0] T389;
  wire[15:0] T253;
  wire[1:0] T254;
  wire[16:0] T255;
  wire[16:0] T256;
  wire[16:0] T257;
  wire[16:0] T390;
  wire[14:0] T258;
  wire[14:0] T391;
  wire[13:0] T259;
  wire[1:0] T260;
  wire[14:0] T261;
  wire[14:0] T262;
  wire[14:0] T263;
  wire[14:0] T392;
  wire[12:0] T264;
  wire[12:0] T393;
  wire[11:0] T265;
  wire[1:0] T266;
  wire[12:0] T267;
  wire[12:0] T268;
  wire[12:0] T269;
  wire[12:0] T394;
  wire[10:0] T270;
  wire[10:0] T395;
  wire[9:0] T271;
  wire[1:0] T272;
  wire[10:0] T273;
  wire[10:0] T274;
  wire[10:0] T275;
  wire[10:0] T396;
  wire[8:0] T276;
  wire[8:0] T397;
  wire[7:0] T277;
  wire[1:0] T278;
  wire[8:0] T279;
  wire[8:0] T280;
  wire[8:0] T281;
  wire[8:0] T398;
  wire[6:0] T282;
  wire[6:0] T399;
  wire[5:0] T283;
  wire[1:0] T284;
  wire[6:0] T285;
  wire[6:0] T286;
  wire[6:0] T287;
  wire[6:0] T400;
  wire[4:0] T288;
  wire[4:0] T401;
  wire[3:0] T289;
  wire[1:0] T290;
  wire[4:0] T291;
  wire[4:0] T292;
  wire[4:0] T293;
  wire[4:0] T402;
  wire[2:0] T294;
  wire[2:0] T403;
  wire[1:0] T295;
  wire[1:0] T296;
  wire[2:0] T297;
  wire[2:0] T298;
  wire[2:0] T299;
  wire[1:0] T300;
  wire[1:0] T301;
  wire[1:0] T302;
  wire[1:0] T303;
  wire[7:0] LogicBlockInBBMuxModule_X_in;


  assign T304 = T0[5'h17:1'h0];
  assign T0 = T3 | T305;
  assign T305 = {1'h0, T1};
  assign T1 = T2 << 5'h12;
  assign T2 = io_config_X_in_3 & 6'h3f;
  assign T3 = T306 & T4;
  assign T4 = ~ T5;
  assign T5 = 25'hfc0000;
  assign T306 = {6'h0, T6};
  assign T6 = T9 | T307;
  assign T307 = {1'h0, T7};
  assign T7 = T8 << 4'hc;
  assign T8 = io_config_X_in_2 & 6'h3f;
  assign T9 = T308 & T10;
  assign T10 = ~ T11;
  assign T11 = 19'h3f000;
  assign T308 = {6'h0, T12};
  assign T12 = T15 | T309;
  assign T309 = {1'h0, T13};
  assign T13 = T14 << 3'h6;
  assign T14 = io_config_X_in_1 & 6'h3f;
  assign T15 = T310 & T16;
  assign T16 = ~ T17;
  assign T17 = 13'hfc0;
  assign T310 = {6'h0, T18};
  assign T18 = T21 | T311;
  assign T311 = {1'h0, T19};
  assign T19 = T20 << 1'h0;
  assign T20 = io_config_X_in_0 & 6'h3f;
  assign T21 = 7'h0 & T22;
  assign T22 = ~ T23;
  assign T23 = 7'h3f;
  assign T312 = T24[3'h7:1'h0];
  assign T24 = T27 | T313;
  assign T313 = {1'h0, T25};
  assign T25 = T26 << 3'h6;
  assign T26 = io_G_wire_below_in_3 & 2'h3;
  assign T27 = T314 & T28;
  assign T28 = ~ T29;
  assign T29 = 9'hc0;
  assign T314 = {2'h0, T30};
  assign T30 = T33 | T315;
  assign T315 = {1'h0, T31};
  assign T31 = T32 << 3'h4;
  assign T32 = io_G_wire_below_in_2 & 2'h3;
  assign T33 = T316 & T34;
  assign T34 = ~ T35;
  assign T35 = 7'h30;
  assign T316 = {2'h0, T36};
  assign T36 = T39 | T317;
  assign T317 = {1'h0, T37};
  assign T37 = T38 << 2'h2;
  assign T38 = io_G_wire_below_in_1 & 2'h3;
  assign T39 = T318 & T40;
  assign T40 = ~ T41;
  assign T41 = 5'hc;
  assign T318 = {2'h0, T42};
  assign T42 = T45 | T319;
  assign T319 = {1'h0, T43};
  assign T43 = T44 << 1'h0;
  assign T44 = io_G_wire_below_in_0 & 2'h3;
  assign T45 = 3'h0 & T46;
  assign T46 = ~ T47;
  assign T47 = 3'h3;
  assign T320 = T48[3'h7:1'h0];
  assign T48 = T51 | T321;
  assign T321 = {1'h0, T49};
  assign T49 = T50 << 3'h6;
  assign T50 = io_G_wire_above_in_3 & 2'h3;
  assign T51 = T322 & T52;
  assign T52 = ~ T53;
  assign T53 = 9'hc0;
  assign T322 = {2'h0, T54};
  assign T54 = T57 | T323;
  assign T323 = {1'h0, T55};
  assign T55 = T56 << 3'h4;
  assign T56 = io_G_wire_above_in_2 & 2'h3;
  assign T57 = T324 & T58;
  assign T58 = ~ T59;
  assign T59 = 7'h30;
  assign T324 = {2'h0, T60};
  assign T60 = T63 | T325;
  assign T325 = {1'h0, T61};
  assign T61 = T62 << 2'h2;
  assign T62 = io_G_wire_above_in_1 & 2'h3;
  assign T63 = T326 & T64;
  assign T64 = ~ T65;
  assign T65 = 5'hc;
  assign T326 = {2'h0, T66};
  assign T66 = T69 | T327;
  assign T327 = {1'h0, T67};
  assign T67 = T68 << 1'h0;
  assign T68 = io_G_wire_above_in_0 & 2'h3;
  assign T69 = 3'h0 & T70;
  assign T70 = ~ T71;
  assign T71 = 3'h3;
  assign T328 = T72[5'h15:1'h0];
  assign T72 = T75 | T329;
  assign T329 = {1'h0, T73};
  assign T73 = T74 << 5'h14;
  assign T74 = io_H_wire_below_in_10 & 2'h3;
  assign T75 = T330 & T76;
  assign T76 = ~ T77;
  assign T77 = 23'h300000;
  assign T330 = {2'h0, T78};
  assign T78 = T81 | T331;
  assign T331 = {1'h0, T79};
  assign T79 = T80 << 5'h12;
  assign T80 = io_H_wire_below_in_9 & 2'h3;
  assign T81 = T332 & T82;
  assign T82 = ~ T83;
  assign T83 = 21'hc0000;
  assign T332 = {2'h0, T84};
  assign T84 = T87 | T333;
  assign T333 = {1'h0, T85};
  assign T85 = T86 << 5'h10;
  assign T86 = io_H_wire_below_in_8 & 2'h3;
  assign T87 = T334 & T88;
  assign T88 = ~ T89;
  assign T89 = 19'h30000;
  assign T334 = {2'h0, T90};
  assign T90 = T93 | T335;
  assign T335 = {1'h0, T91};
  assign T91 = T92 << 4'he;
  assign T92 = io_H_wire_below_in_7 & 2'h3;
  assign T93 = T336 & T94;
  assign T94 = ~ T95;
  assign T95 = 17'hc000;
  assign T336 = {2'h0, T96};
  assign T96 = T99 | T337;
  assign T337 = {1'h0, T97};
  assign T97 = T98 << 4'hc;
  assign T98 = io_H_wire_below_in_6 & 2'h3;
  assign T99 = T338 & T100;
  assign T100 = ~ T101;
  assign T101 = 15'h3000;
  assign T338 = {2'h0, T102};
  assign T102 = T105 | T339;
  assign T339 = {1'h0, T103};
  assign T103 = T104 << 4'ha;
  assign T104 = io_H_wire_below_in_5 & 2'h3;
  assign T105 = T340 & T106;
  assign T106 = ~ T107;
  assign T107 = 13'hc00;
  assign T340 = {2'h0, T108};
  assign T108 = T111 | T341;
  assign T341 = {1'h0, T109};
  assign T109 = T110 << 4'h8;
  assign T110 = io_H_wire_below_in_4 & 2'h3;
  assign T111 = T342 & T112;
  assign T112 = ~ T113;
  assign T113 = 11'h300;
  assign T342 = {2'h0, T114};
  assign T114 = T117 | T343;
  assign T343 = {1'h0, T115};
  assign T115 = T116 << 3'h6;
  assign T116 = io_H_wire_below_in_3 & 2'h3;
  assign T117 = T344 & T118;
  assign T118 = ~ T119;
  assign T119 = 9'hc0;
  assign T344 = {2'h0, T120};
  assign T120 = T123 | T345;
  assign T345 = {1'h0, T121};
  assign T121 = T122 << 3'h4;
  assign T122 = io_H_wire_below_in_2 & 2'h3;
  assign T123 = T346 & T124;
  assign T124 = ~ T125;
  assign T125 = 7'h30;
  assign T346 = {2'h0, T126};
  assign T126 = T129 | T347;
  assign T347 = {1'h0, T127};
  assign T127 = T128 << 2'h2;
  assign T128 = io_H_wire_below_in_1 & 2'h3;
  assign T129 = T348 & T130;
  assign T130 = ~ T131;
  assign T131 = 5'hc;
  assign T348 = {2'h0, T132};
  assign T132 = T135 | T349;
  assign T349 = {1'h0, T133};
  assign T133 = T134 << 1'h0;
  assign T134 = io_H_wire_below_in_0 & 2'h3;
  assign T135 = 3'h0 & T136;
  assign T136 = ~ T137;
  assign T137 = 3'h3;
  assign T350 = T138[5'h15:1'h0];
  assign T138 = T141 | T351;
  assign T351 = {1'h0, T139};
  assign T139 = T140 << 5'h14;
  assign T140 = io_H_wire_above_in_10 & 2'h3;
  assign T141 = T352 & T142;
  assign T142 = ~ T143;
  assign T143 = 23'h300000;
  assign T352 = {2'h0, T144};
  assign T144 = T147 | T353;
  assign T353 = {1'h0, T145};
  assign T145 = T146 << 5'h12;
  assign T146 = io_H_wire_above_in_9 & 2'h3;
  assign T147 = T354 & T148;
  assign T148 = ~ T149;
  assign T149 = 21'hc0000;
  assign T354 = {2'h0, T150};
  assign T150 = T153 | T355;
  assign T355 = {1'h0, T151};
  assign T151 = T152 << 5'h10;
  assign T152 = io_H_wire_above_in_8 & 2'h3;
  assign T153 = T356 & T154;
  assign T154 = ~ T155;
  assign T155 = 19'h30000;
  assign T356 = {2'h0, T156};
  assign T156 = T159 | T357;
  assign T357 = {1'h0, T157};
  assign T157 = T158 << 4'he;
  assign T158 = io_H_wire_above_in_7 & 2'h3;
  assign T159 = T358 & T160;
  assign T160 = ~ T161;
  assign T161 = 17'hc000;
  assign T358 = {2'h0, T162};
  assign T162 = T165 | T359;
  assign T359 = {1'h0, T163};
  assign T163 = T164 << 4'hc;
  assign T164 = io_H_wire_above_in_6 & 2'h3;
  assign T165 = T360 & T166;
  assign T166 = ~ T167;
  assign T167 = 15'h3000;
  assign T360 = {2'h0, T168};
  assign T168 = T171 | T361;
  assign T361 = {1'h0, T169};
  assign T169 = T170 << 4'ha;
  assign T170 = io_H_wire_above_in_5 & 2'h3;
  assign T171 = T362 & T172;
  assign T172 = ~ T173;
  assign T173 = 13'hc00;
  assign T362 = {2'h0, T174};
  assign T174 = T177 | T363;
  assign T363 = {1'h0, T175};
  assign T175 = T176 << 4'h8;
  assign T176 = io_H_wire_above_in_4 & 2'h3;
  assign T177 = T364 & T178;
  assign T178 = ~ T179;
  assign T179 = 11'h300;
  assign T364 = {2'h0, T180};
  assign T180 = T183 | T365;
  assign T365 = {1'h0, T181};
  assign T181 = T182 << 3'h6;
  assign T182 = io_H_wire_above_in_3 & 2'h3;
  assign T183 = T366 & T184;
  assign T184 = ~ T185;
  assign T185 = 9'hc0;
  assign T366 = {2'h0, T186};
  assign T186 = T189 | T367;
  assign T367 = {1'h0, T187};
  assign T187 = T188 << 3'h4;
  assign T188 = io_H_wire_above_in_2 & 2'h3;
  assign T189 = T368 & T190;
  assign T190 = ~ T191;
  assign T191 = 7'h30;
  assign T368 = {2'h0, T192};
  assign T192 = T195 | T369;
  assign T369 = {1'h0, T193};
  assign T193 = T194 << 2'h2;
  assign T194 = io_H_wire_above_in_1 & 2'h3;
  assign T195 = T370 & T196;
  assign T196 = ~ T197;
  assign T197 = 5'hc;
  assign T370 = {2'h0, T198};
  assign T198 = T201 | T371;
  assign T371 = {1'h0, T199};
  assign T199 = T200 << 1'h0;
  assign T200 = io_H_wire_above_in_0 & 2'h3;
  assign T201 = 3'h0 & T202;
  assign T202 = ~ T203;
  assign T203 = 3'h3;
  assign T372 = T204[5'h1f:1'h0];
  assign T204 = T207 | T373;
  assign T373 = {1'h0, T205};
  assign T205 = T206 << 5'h1e;
  assign T206 = io_V_wire_in_15 & 2'h3;
  assign T207 = T374 & T208;
  assign T208 = ~ T209;
  assign T209 = 33'hc0000000;
  assign T374 = {2'h0, T210};
  assign T210 = T213 | T375;
  assign T375 = {1'h0, T211};
  assign T211 = T212 << 5'h1c;
  assign T212 = io_V_wire_in_14 & 2'h3;
  assign T213 = T376 & T214;
  assign T214 = ~ T215;
  assign T215 = 31'h30000000;
  assign T376 = {2'h0, T216};
  assign T216 = T219 | T377;
  assign T377 = {1'h0, T217};
  assign T217 = T218 << 5'h1a;
  assign T218 = io_V_wire_in_13 & 2'h3;
  assign T219 = T378 & T220;
  assign T220 = ~ T221;
  assign T221 = 29'hc000000;
  assign T378 = {2'h0, T222};
  assign T222 = T225 | T379;
  assign T379 = {1'h0, T223};
  assign T223 = T224 << 5'h18;
  assign T224 = io_V_wire_in_12 & 2'h3;
  assign T225 = T380 & T226;
  assign T226 = ~ T227;
  assign T227 = 27'h3000000;
  assign T380 = {2'h0, T228};
  assign T228 = T231 | T381;
  assign T381 = {1'h0, T229};
  assign T229 = T230 << 5'h16;
  assign T230 = io_V_wire_in_11 & 2'h3;
  assign T231 = T382 & T232;
  assign T232 = ~ T233;
  assign T233 = 25'hc00000;
  assign T382 = {2'h0, T234};
  assign T234 = T237 | T383;
  assign T383 = {1'h0, T235};
  assign T235 = T236 << 5'h14;
  assign T236 = io_V_wire_in_10 & 2'h3;
  assign T237 = T384 & T238;
  assign T238 = ~ T239;
  assign T239 = 23'h300000;
  assign T384 = {2'h0, T240};
  assign T240 = T243 | T385;
  assign T385 = {1'h0, T241};
  assign T241 = T242 << 5'h12;
  assign T242 = io_V_wire_in_9 & 2'h3;
  assign T243 = T386 & T244;
  assign T244 = ~ T245;
  assign T245 = 21'hc0000;
  assign T386 = {2'h0, T246};
  assign T246 = T249 | T387;
  assign T387 = {1'h0, T247};
  assign T247 = T248 << 5'h10;
  assign T248 = io_V_wire_in_8 & 2'h3;
  assign T249 = T388 & T250;
  assign T250 = ~ T251;
  assign T251 = 19'h30000;
  assign T388 = {2'h0, T252};
  assign T252 = T255 | T389;
  assign T389 = {1'h0, T253};
  assign T253 = T254 << 4'he;
  assign T254 = io_V_wire_in_7 & 2'h3;
  assign T255 = T390 & T256;
  assign T256 = ~ T257;
  assign T257 = 17'hc000;
  assign T390 = {2'h0, T258};
  assign T258 = T261 | T391;
  assign T391 = {1'h0, T259};
  assign T259 = T260 << 4'hc;
  assign T260 = io_V_wire_in_6 & 2'h3;
  assign T261 = T392 & T262;
  assign T262 = ~ T263;
  assign T263 = 15'h3000;
  assign T392 = {2'h0, T264};
  assign T264 = T267 | T393;
  assign T393 = {1'h0, T265};
  assign T265 = T266 << 4'ha;
  assign T266 = io_V_wire_in_5 & 2'h3;
  assign T267 = T394 & T268;
  assign T268 = ~ T269;
  assign T269 = 13'hc00;
  assign T394 = {2'h0, T270};
  assign T270 = T273 | T395;
  assign T395 = {1'h0, T271};
  assign T271 = T272 << 4'h8;
  assign T272 = io_V_wire_in_4 & 2'h3;
  assign T273 = T396 & T274;
  assign T274 = ~ T275;
  assign T275 = 11'h300;
  assign T396 = {2'h0, T276};
  assign T276 = T279 | T397;
  assign T397 = {1'h0, T277};
  assign T277 = T278 << 3'h6;
  assign T278 = io_V_wire_in_3 & 2'h3;
  assign T279 = T398 & T280;
  assign T280 = ~ T281;
  assign T281 = 9'hc0;
  assign T398 = {2'h0, T282};
  assign T282 = T285 | T399;
  assign T399 = {1'h0, T283};
  assign T283 = T284 << 3'h4;
  assign T284 = io_V_wire_in_2 & 2'h3;
  assign T285 = T400 & T286;
  assign T286 = ~ T287;
  assign T287 = 7'h30;
  assign T400 = {2'h0, T288};
  assign T288 = T291 | T401;
  assign T401 = {1'h0, T289};
  assign T289 = T290 << 2'h2;
  assign T290 = io_V_wire_in_1 & 2'h3;
  assign T291 = T402 & T292;
  assign T292 = ~ T293;
  assign T293 = 5'hc;
  assign T402 = {2'h0, T294};
  assign T294 = T297 | T403;
  assign T403 = {1'h0, T295};
  assign T295 = T296 << 1'h0;
  assign T296 = io_V_wire_in_0 & 2'h3;
  assign T297 = 3'h0 & T298;
  assign T298 = ~ T299;
  assign T299 = 3'h3;
  assign io_X_in_0 = T300;
  assign T300 = LogicBlockInBBMuxModule_X_in[1'h1:1'h0];
  assign io_X_in_1 = T301;
  assign T301 = LogicBlockInBBMuxModule_X_in[2'h3:2'h2];
  assign io_X_in_2 = T302;
  assign T302 = LogicBlockInBBMuxModule_X_in[3'h5:3'h4];
  assign io_X_in_3 = T303;
  assign T303 = LogicBlockInBBMuxModule_X_in[3'h7:3'h6];
  input_mux LogicBlockInBBMuxModule(
       .V_wire_in( T372 ),
       .H_wire_above_in( T350 ),
       .H_wire_below_in( T328 ),
       .G_wire_above_in( T320 ),
       .G_wire_below_in( T312 ),
       .config_X_in( T304 ),
       .Z_reg( io_Z_reg ),
       .D_reg( io_D_reg ),
       .X_in( LogicBlockInBBMuxModule_X_in )
  );
endmodule

module CrossbarModule(
    input [1:0] io_in,
    input [1:0] io_sel,
    output[1:0] io_out
);

  wire[1:0] T42;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T43;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire[1:0] T44;
  wire T7;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire[1:0] T45;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[2:0] T46;
  wire T26;
  wire T27;
  wire T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T47;
  wire T31;
  wire T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire[2:0] T48;
  wire T36;
  wire T37;
  wire T38;
  wire[2:0] T39;
  wire[2:0] T40;
  wire T41;


  assign io_out = T42;
  assign T42 = T0[1'h1:1'h0];
  assign T0 = T41 ? T33 : T1;
  assign T1 = T31 ? T23 : T43;
  assign T43 = {1'h0, T2};
  assign T2 = T22 ? T14 : T3;
  assign T3 = T12 ? T4 : 2'h0;
  assign T4 = T10 | T5;
  assign T5 = T44 & T6;
  assign T6 = 2'h1;
  assign T44 = T7 ? 2'h3 : 2'h0;
  assign T7 = T8;
  assign T8 = T9;
  assign T9 = io_in[1'h0];
  assign T10 = 2'h0 & T11;
  assign T11 = ~ T6;
  assign T12 = T13 == 1'h0;
  assign T13 = io_sel[1'h0];
  assign T14 = T20 | T15;
  assign T15 = T45 & T16;
  assign T16 = 2'h1;
  assign T45 = T17 ? 2'h3 : 2'h0;
  assign T17 = T18;
  assign T18 = T19;
  assign T19 = io_in[1'h1];
  assign T20 = T3 & T21;
  assign T21 = ~ T16;
  assign T22 = T12 ^ 1'h1;
  assign T23 = T29 | T24;
  assign T24 = T46 & T25;
  assign T25 = 3'h2;
  assign T46 = T26 ? 3'h7 : 3'h0;
  assign T26 = T27;
  assign T27 = T28;
  assign T28 = io_in[1'h0];
  assign T29 = T47 & T30;
  assign T30 = ~ T25;
  assign T47 = {1'h0, T2};
  assign T31 = T32 == 1'h0;
  assign T32 = io_sel[1'h1];
  assign T33 = T39 | T34;
  assign T34 = T48 & T35;
  assign T35 = 3'h2;
  assign T48 = T36 ? 3'h7 : 3'h0;
  assign T36 = T37;
  assign T37 = T38;
  assign T38 = io_in[1'h1];
  assign T39 = T1 & T40;
  assign T40 = ~ T35;
  assign T41 = T31 ^ 1'h1;
endmodule

module ShiftInvertModule(
    input  io_shift_in,
    input [1:0] io_in,
    input [1:0] io_sel,
    output[1:0] io_out,
    output io_shift_out
);

  wire T0;
  wire[1:0] T80;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T81;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T82;
  wire T12;
  wire T13;
  wire T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T83;
  wire T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T84;
  wire T25;
  wire[2:0] T26;
  wire[2:0] T85;
  wire[1:0] T27;
  wire[1:0] T28;
  wire[1:0] T86;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T87;
  wire[2:0] T33;
  wire[2:0] T88;
  wire[1:0] T34;
  wire T89;
  wire[2:0] T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire[2:0] T90;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire[2:0] T42;
  wire[2:0] T43;
  wire T44;
  wire[2:0] T45;
  wire[2:0] T91;
  wire[1:0] T46;
  wire[1:0] T47;
  wire[1:0] T92;
  wire T48;
  wire T49;
  wire T93;
  wire[2:0] T50;
  wire[2:0] T94;
  wire[1:0] T51;
  wire T95;
  wire[2:0] T52;
  wire[2:0] T53;
  wire[2:0] T54;
  wire[2:0] T96;
  wire T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire[2:0] T59;
  wire T60;
  wire[2:0] T61;
  wire[2:0] T97;
  wire[1:0] T62;
  wire[1:0] T63;
  wire[1:0] T98;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T99;
  wire[2:0] T68;
  wire[2:0] T100;
  wire[1:0] T69;
  wire T101;
  wire[2:0] T70;
  wire[2:0] T71;
  wire[2:0] T72;
  wire[2:0] T102;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[2:0] T77;
  wire[2:0] T78;
  wire T79;


  assign io_shift_out = T0;
  assign T0 = io_in[1'h1];
  assign io_out = T80;
  assign T80 = T1[1'h1:1'h0];
  assign T1 = T79 ? T70 : T2;
  assign T2 = T79 ? T61 : T3;
  assign T3 = T60 ? T52 : T4;
  assign T4 = T60 ? T45 : T5;
  assign T5 = T44 ? T35 : T6;
  assign T6 = T44 ? T26 : T7;
  assign T7 = T25 ? T17 : T81;
  assign T81 = {1'h0, T8};
  assign T8 = T25 ? T9 : 2'h0;
  assign T9 = T15 | T10;
  assign T10 = T82 & T11;
  assign T11 = 2'h1;
  assign T82 = T12 ? 2'h3 : 2'h0;
  assign T12 = T13;
  assign T13 = T14;
  assign T14 = io_in[1'h0];
  assign T15 = 2'h0 & T16;
  assign T16 = ~ T11;
  assign T17 = T23 | T18;
  assign T18 = T83 & T19;
  assign T19 = 3'h2;
  assign T83 = T20 ? 3'h7 : 3'h0;
  assign T20 = T21;
  assign T21 = T22;
  assign T22 = io_in[1'h1];
  assign T23 = T84 & T24;
  assign T24 = ~ T19;
  assign T84 = {1'h0, T8};
  assign T25 = 2'h0 == io_sel;
  assign T26 = T33 | T85;
  assign T85 = {T87, T27};
  assign T27 = T86 & T28;
  assign T28 = 2'h1;
  assign T86 = T29 ? 2'h3 : 2'h0;
  assign T29 = T30;
  assign T30 = T31;
  assign T31 = ~ T32;
  assign T32 = io_in[1'h0];
  assign T87 = T27[1'h1];
  assign T33 = T7 & T88;
  assign T88 = {T89, T34};
  assign T34 = ~ T28;
  assign T89 = T34[1'h1];
  assign T35 = T42 | T36;
  assign T36 = T90 & T37;
  assign T37 = 3'h2;
  assign T90 = T38 ? 3'h7 : 3'h0;
  assign T38 = T39;
  assign T39 = T40;
  assign T40 = ~ T41;
  assign T41 = io_in[1'h1];
  assign T42 = T6 & T43;
  assign T43 = ~ T37;
  assign T44 = 2'h1 == io_sel;
  assign T45 = T50 | T91;
  assign T91 = {T93, T46};
  assign T46 = T92 & T47;
  assign T47 = 2'h1;
  assign T92 = T48 ? 2'h3 : 2'h0;
  assign T48 = T49;
  assign T49 = io_shift_in;
  assign T93 = T46[1'h1];
  assign T50 = T5 & T94;
  assign T94 = {T95, T51};
  assign T51 = ~ T47;
  assign T95 = T51[1'h1];
  assign T52 = T58 | T53;
  assign T53 = T96 & T54;
  assign T54 = 3'h2;
  assign T96 = T55 ? 3'h7 : 3'h0;
  assign T55 = T56;
  assign T56 = T57;
  assign T57 = io_in[1'h0];
  assign T58 = T4 & T59;
  assign T59 = ~ T54;
  assign T60 = 2'h2 == io_sel;
  assign T61 = T68 | T97;
  assign T97 = {T99, T62};
  assign T62 = T98 & T63;
  assign T63 = 2'h1;
  assign T98 = T64 ? 2'h3 : 2'h0;
  assign T64 = T65;
  assign T65 = T66;
  assign T66 = T67;
  assign T67 = ~ io_shift_in;
  assign T99 = T62[1'h1];
  assign T68 = T3 & T100;
  assign T100 = {T101, T69};
  assign T69 = ~ T63;
  assign T101 = T69[1'h1];
  assign T70 = T77 | T71;
  assign T71 = T102 & T72;
  assign T72 = 3'h2;
  assign T102 = T73 ? 3'h7 : 3'h0;
  assign T73 = T74;
  assign T74 = T75;
  assign T75 = ~ T76;
  assign T76 = io_in[1'h0];
  assign T77 = T2 & T78;
  assign T78 = ~ T72;
  assign T79 = 2'h3 == io_sel;
endmodule

module CarrySaveAdderModule(
    input  io_shift_carry_in,
    input [1:0] io_in_2,
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    output[1:0] io_sum,
    output[1:0] io_carry,
    output io_shift_carry_out
);

  wire T0;
  wire[1:0] carry;
  wire[1:0] T76;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T77;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T78;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[1:0] T79;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T80;
  wire[2:0] T37;
  wire[2:0] T81;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T82;
  wire T40;
  wire T41;
  wire T83;
  wire[2:0] T42;
  wire[2:0] T84;
  wire[1:0] T43;
  wire T85;
  wire[2:0] T44;
  wire[2:0] T45;
  wire[2:0] T46;
  wire[2:0] T86;
  wire T47;
  wire T48;
  wire T49;
  wire[2:0] T50;
  wire[2:0] T51;
  wire[1:0] T87;
  wire[2:0] T52;
  wire[2:0] T53;
  wire[2:0] T54;
  wire[2:0] T88;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[2:0] T63;
  wire[2:0] T89;
  wire[1:0] T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T90;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire[1:0] T74;
  wire[1:0] T75;


  assign io_shift_carry_out = T0;
  assign T0 = carry[1'h1];
  assign carry = T76;
  assign T76 = T1[1'h1:1'h0];
  assign T1 = T17 | T2;
  assign T2 = T77 & T3;
  assign T3 = 3'h2;
  assign T77 = T4 ? 3'h7 : 3'h0;
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = T10 | T7;
  assign T7 = T9 & T8;
  assign T8 = io_in_0[1'h1];
  assign T9 = io_in_2[1'h1];
  assign T10 = T14 | T11;
  assign T11 = T13 & T12;
  assign T12 = io_in_0[1'h1];
  assign T13 = io_in_1[1'h1];
  assign T14 = T16 & T15;
  assign T15 = io_in_1[1'h1];
  assign T16 = io_in_2[1'h1];
  assign T17 = T78 & T18;
  assign T18 = ~ T3;
  assign T78 = {1'h0, T19};
  assign T19 = T35 | T20;
  assign T20 = T79 & T21;
  assign T21 = 2'h1;
  assign T79 = T22 ? 2'h3 : 2'h0;
  assign T22 = T23;
  assign T23 = T24;
  assign T24 = T28 | T25;
  assign T25 = T27 & T26;
  assign T26 = io_in_0[1'h0];
  assign T27 = io_in_2[1'h0];
  assign T28 = T32 | T29;
  assign T29 = T31 & T30;
  assign T30 = io_in_0[1'h0];
  assign T31 = io_in_1[1'h0];
  assign T32 = T34 & T33;
  assign T33 = io_in_1[1'h0];
  assign T34 = io_in_2[1'h0];
  assign T35 = 2'h0 & T36;
  assign T36 = ~ T21;
  assign io_carry = T80;
  assign T80 = T37[1'h1:1'h0];
  assign T37 = T42 | T81;
  assign T81 = {T83, T38};
  assign T38 = T82 & T39;
  assign T39 = 2'h1;
  assign T82 = T40 ? 2'h3 : 2'h0;
  assign T40 = T41;
  assign T41 = io_shift_carry_in;
  assign T83 = T38[1'h1];
  assign T42 = T44 & T84;
  assign T84 = {T85, T43};
  assign T43 = ~ T39;
  assign T85 = T43[1'h1];
  assign T44 = T50 | T45;
  assign T45 = T86 & T46;
  assign T46 = 3'h2;
  assign T86 = T47 ? 3'h7 : 3'h0;
  assign T47 = T48;
  assign T48 = T49;
  assign T49 = carry[1'h0];
  assign T50 = 3'h0 & T51;
  assign T51 = ~ T46;
  assign io_sum = T87;
  assign T87 = T52[1'h1:1'h0];
  assign T52 = T62 | T53;
  assign T53 = T88 & T54;
  assign T54 = 3'h2;
  assign T88 = T55 ? 3'h7 : 3'h0;
  assign T55 = T56;
  assign T56 = T57;
  assign T57 = T59 ^ T58;
  assign T58 = io_in_0[1'h1];
  assign T59 = T61 ^ T60;
  assign T60 = io_in_1[1'h1];
  assign T61 = io_in_2[1'h1];
  assign T62 = T89 & T63;
  assign T63 = ~ T54;
  assign T89 = {1'h0, T64};
  assign T64 = T74 | T65;
  assign T65 = T90 & T66;
  assign T66 = 2'h1;
  assign T90 = T67 ? 2'h3 : 2'h0;
  assign T67 = T68;
  assign T68 = T69;
  assign T69 = T71 ^ T70;
  assign T70 = io_in_0[1'h0];
  assign T71 = T73 ^ T72;
  assign T72 = io_in_1[1'h0];
  assign T73 = io_in_2[1'h0];
  assign T74 = 2'h0 & T75;
  assign T75 = ~ T66;
endmodule

module LookUpTableModule(
    input [1:0] io_in_2,
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    input [7:0] io_config,
    output[1:0] io_out
);

  wire[1:0] T208;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T209;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire[1:0] T210;
  wire T19;
  wire T20;
  wire T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire T24;
  wire[2:0] in_0;
  wire[2:0] T211;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] T212;
  wire T28;
  wire T29;
  wire T30;
  wire[3:0] T31;
  wire[3:0] T32;
  wire[3:0] T213;
  wire[2:0] T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire[2:0] T214;
  wire T36;
  wire T37;
  wire T38;
  wire[2:0] T39;
  wire[2:0] T40;
  wire[2:0] T215;
  wire[1:0] T41;
  wire[1:0] T42;
  wire[1:0] T43;
  wire[1:0] T216;
  wire T44;
  wire T45;
  wire T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire[1:0] T50;
  wire[1:0] T51;
  wire[1:0] T217;
  wire T52;
  wire T53;
  wire T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire[1:0] T60;
  wire[1:0] T218;
  wire T61;
  wire T62;
  wire T63;
  wire[1:0] T64;
  wire[1:0] T65;
  wire T66;
  wire[1:0] T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire[1:0] T219;
  wire T70;
  wire T71;
  wire T72;
  wire[1:0] T73;
  wire[1:0] T74;
  wire T75;
  wire[1:0] T76;
  wire[1:0] T77;
  wire[1:0] T78;
  wire[1:0] T220;
  wire T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire[1:0] T83;
  wire T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire[1:0] T221;
  wire T88;
  wire T89;
  wire T90;
  wire[1:0] T91;
  wire[1:0] T92;
  wire T93;
  wire[1:0] T94;
  wire[1:0] T95;
  wire[1:0] T96;
  wire[1:0] T222;
  wire T97;
  wire T98;
  wire T99;
  wire[1:0] T100;
  wire[1:0] T101;
  wire T102;
  wire[1:0] T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire[1:0] T223;
  wire T106;
  wire T107;
  wire T108;
  wire[1:0] T109;
  wire[1:0] T110;
  wire T111;
  wire[2:0] T112;
  wire[2:0] T113;
  wire[2:0] T114;
  wire[2:0] T224;
  wire T115;
  wire T116;
  wire T117;
  wire[2:0] T118;
  wire[2:0] T119;
  wire[2:0] T225;
  wire T120;
  wire[2:0] in_1;
  wire[2:0] T226;
  wire[3:0] T121;
  wire[3:0] T122;
  wire[3:0] T123;
  wire[3:0] T227;
  wire T124;
  wire T125;
  wire T126;
  wire[3:0] T127;
  wire[3:0] T128;
  wire[3:0] T228;
  wire[2:0] T129;
  wire[2:0] T130;
  wire[2:0] T131;
  wire[2:0] T229;
  wire T132;
  wire T133;
  wire T134;
  wire[2:0] T135;
  wire[2:0] T136;
  wire[2:0] T230;
  wire[1:0] T137;
  wire[1:0] T138;
  wire[1:0] T139;
  wire[1:0] T231;
  wire T140;
  wire T141;
  wire T142;
  wire[1:0] T143;
  wire[1:0] T144;
  wire[2:0] T145;
  wire[2:0] T146;
  wire[2:0] T147;
  wire[2:0] T232;
  wire T148;
  wire T149;
  wire T150;
  wire[2:0] T151;
  wire[2:0] T152;
  wire T153;
  wire[2:0] T154;
  wire[2:0] T155;
  wire[2:0] T156;
  wire[2:0] T233;
  wire T157;
  wire T158;
  wire T159;
  wire[2:0] T160;
  wire[2:0] T161;
  wire T162;
  wire[2:0] T163;
  wire[2:0] T164;
  wire[2:0] T165;
  wire[2:0] T234;
  wire T166;
  wire T167;
  wire T168;
  wire[2:0] T169;
  wire[2:0] T170;
  wire T171;
  wire[2:0] T172;
  wire[2:0] T173;
  wire[2:0] T174;
  wire[2:0] T235;
  wire T175;
  wire T176;
  wire T177;
  wire[2:0] T178;
  wire[2:0] T179;
  wire T180;
  wire[2:0] T181;
  wire[2:0] T182;
  wire[2:0] T183;
  wire[2:0] T236;
  wire T184;
  wire T185;
  wire T186;
  wire[2:0] T187;
  wire[2:0] T188;
  wire T189;
  wire[2:0] T190;
  wire[2:0] T191;
  wire[2:0] T192;
  wire[2:0] T237;
  wire T193;
  wire T194;
  wire T195;
  wire[2:0] T196;
  wire[2:0] T197;
  wire T198;
  wire[2:0] T199;
  wire[2:0] T200;
  wire[2:0] T201;
  wire[2:0] T238;
  wire T202;
  wire T203;
  wire T204;
  wire[2:0] T205;
  wire[2:0] T206;
  wire T207;


  assign io_out = T208;
  assign T208 = T0[1'h1:1'h0];
  assign T0 = T207 ? T199 : T1;
  assign T1 = T198 ? T190 : T2;
  assign T2 = T189 ? T181 : T3;
  assign T3 = T180 ? T172 : T4;
  assign T4 = T171 ? T163 : T5;
  assign T5 = T162 ? T154 : T6;
  assign T6 = T153 ? T145 : T7;
  assign T7 = T120 ? T112 : T209;
  assign T209 = {1'h0, T8};
  assign T8 = T111 ? T103 : T9;
  assign T9 = T102 ? T94 : T10;
  assign T10 = T93 ? T85 : T11;
  assign T11 = T84 ? T76 : T12;
  assign T12 = T75 ? T67 : T13;
  assign T13 = T66 ? T58 : T14;
  assign T14 = T57 ? T49 : T15;
  assign T15 = T24 ? T16 : 2'h0;
  assign T16 = T22 | T17;
  assign T17 = T210 & T18;
  assign T18 = 2'h1;
  assign T210 = T19 ? 2'h3 : 2'h0;
  assign T19 = T20;
  assign T20 = T21;
  assign T21 = io_config[1'h0];
  assign T22 = 2'h0 & T23;
  assign T23 = ~ T18;
  assign T24 = 3'h0 == in_0;
  assign in_0 = T211;
  assign T211 = T25[2'h2:1'h0];
  assign T25 = T31 | T26;
  assign T26 = T212 & T27;
  assign T27 = 4'h4;
  assign T212 = T28 ? 4'hf : 4'h0;
  assign T28 = T29;
  assign T29 = T30;
  assign T30 = io_in_2[1'h0];
  assign T31 = T213 & T32;
  assign T32 = ~ T27;
  assign T213 = {1'h0, T33};
  assign T33 = T39 | T34;
  assign T34 = T214 & T35;
  assign T35 = 3'h2;
  assign T214 = T36 ? 3'h7 : 3'h0;
  assign T36 = T37;
  assign T37 = T38;
  assign T38 = io_in_1[1'h0];
  assign T39 = T215 & T40;
  assign T40 = ~ T35;
  assign T215 = {1'h0, T41};
  assign T41 = T47 | T42;
  assign T42 = T216 & T43;
  assign T43 = 2'h1;
  assign T216 = T44 ? 2'h3 : 2'h0;
  assign T44 = T45;
  assign T45 = T46;
  assign T46 = io_in_0[1'h0];
  assign T47 = 2'h0 & T48;
  assign T48 = ~ T43;
  assign T49 = T55 | T50;
  assign T50 = T217 & T51;
  assign T51 = 2'h1;
  assign T217 = T52 ? 2'h3 : 2'h0;
  assign T52 = T53;
  assign T53 = T54;
  assign T54 = io_config[1'h1];
  assign T55 = T15 & T56;
  assign T56 = ~ T51;
  assign T57 = 3'h1 == in_0;
  assign T58 = T64 | T59;
  assign T59 = T218 & T60;
  assign T60 = 2'h1;
  assign T218 = T61 ? 2'h3 : 2'h0;
  assign T61 = T62;
  assign T62 = T63;
  assign T63 = io_config[2'h2];
  assign T64 = T14 & T65;
  assign T65 = ~ T60;
  assign T66 = 3'h2 == in_0;
  assign T67 = T73 | T68;
  assign T68 = T219 & T69;
  assign T69 = 2'h1;
  assign T219 = T70 ? 2'h3 : 2'h0;
  assign T70 = T71;
  assign T71 = T72;
  assign T72 = io_config[2'h3];
  assign T73 = T13 & T74;
  assign T74 = ~ T69;
  assign T75 = 3'h3 == in_0;
  assign T76 = T82 | T77;
  assign T77 = T220 & T78;
  assign T78 = 2'h1;
  assign T220 = T79 ? 2'h3 : 2'h0;
  assign T79 = T80;
  assign T80 = T81;
  assign T81 = io_config[3'h4];
  assign T82 = T12 & T83;
  assign T83 = ~ T78;
  assign T84 = 3'h4 == in_0;
  assign T85 = T91 | T86;
  assign T86 = T221 & T87;
  assign T87 = 2'h1;
  assign T221 = T88 ? 2'h3 : 2'h0;
  assign T88 = T89;
  assign T89 = T90;
  assign T90 = io_config[3'h5];
  assign T91 = T11 & T92;
  assign T92 = ~ T87;
  assign T93 = 3'h5 == in_0;
  assign T94 = T100 | T95;
  assign T95 = T222 & T96;
  assign T96 = 2'h1;
  assign T222 = T97 ? 2'h3 : 2'h0;
  assign T97 = T98;
  assign T98 = T99;
  assign T99 = io_config[3'h6];
  assign T100 = T10 & T101;
  assign T101 = ~ T96;
  assign T102 = 3'h6 == in_0;
  assign T103 = T109 | T104;
  assign T104 = T223 & T105;
  assign T105 = 2'h1;
  assign T223 = T106 ? 2'h3 : 2'h0;
  assign T106 = T107;
  assign T107 = T108;
  assign T108 = io_config[3'h7];
  assign T109 = T9 & T110;
  assign T110 = ~ T105;
  assign T111 = 3'h7 == in_0;
  assign T112 = T118 | T113;
  assign T113 = T224 & T114;
  assign T114 = 3'h2;
  assign T224 = T115 ? 3'h7 : 3'h0;
  assign T115 = T116;
  assign T116 = T117;
  assign T117 = io_config[1'h0];
  assign T118 = T225 & T119;
  assign T119 = ~ T114;
  assign T225 = {1'h0, T8};
  assign T120 = 3'h0 == in_1;
  assign in_1 = T226;
  assign T226 = T121[2'h2:1'h0];
  assign T121 = T127 | T122;
  assign T122 = T227 & T123;
  assign T123 = 4'h4;
  assign T227 = T124 ? 4'hf : 4'h0;
  assign T124 = T125;
  assign T125 = T126;
  assign T126 = io_in_2[1'h1];
  assign T127 = T228 & T128;
  assign T128 = ~ T123;
  assign T228 = {1'h0, T129};
  assign T129 = T135 | T130;
  assign T130 = T229 & T131;
  assign T131 = 3'h2;
  assign T229 = T132 ? 3'h7 : 3'h0;
  assign T132 = T133;
  assign T133 = T134;
  assign T134 = io_in_1[1'h1];
  assign T135 = T230 & T136;
  assign T136 = ~ T131;
  assign T230 = {1'h0, T137};
  assign T137 = T143 | T138;
  assign T138 = T231 & T139;
  assign T139 = 2'h1;
  assign T231 = T140 ? 2'h3 : 2'h0;
  assign T140 = T141;
  assign T141 = T142;
  assign T142 = io_in_0[1'h1];
  assign T143 = 2'h0 & T144;
  assign T144 = ~ T139;
  assign T145 = T151 | T146;
  assign T146 = T232 & T147;
  assign T147 = 3'h2;
  assign T232 = T148 ? 3'h7 : 3'h0;
  assign T148 = T149;
  assign T149 = T150;
  assign T150 = io_config[1'h1];
  assign T151 = T7 & T152;
  assign T152 = ~ T147;
  assign T153 = 3'h1 == in_1;
  assign T154 = T160 | T155;
  assign T155 = T233 & T156;
  assign T156 = 3'h2;
  assign T233 = T157 ? 3'h7 : 3'h0;
  assign T157 = T158;
  assign T158 = T159;
  assign T159 = io_config[2'h2];
  assign T160 = T6 & T161;
  assign T161 = ~ T156;
  assign T162 = 3'h2 == in_1;
  assign T163 = T169 | T164;
  assign T164 = T234 & T165;
  assign T165 = 3'h2;
  assign T234 = T166 ? 3'h7 : 3'h0;
  assign T166 = T167;
  assign T167 = T168;
  assign T168 = io_config[2'h3];
  assign T169 = T5 & T170;
  assign T170 = ~ T165;
  assign T171 = 3'h3 == in_1;
  assign T172 = T178 | T173;
  assign T173 = T235 & T174;
  assign T174 = 3'h2;
  assign T235 = T175 ? 3'h7 : 3'h0;
  assign T175 = T176;
  assign T176 = T177;
  assign T177 = io_config[3'h4];
  assign T178 = T4 & T179;
  assign T179 = ~ T174;
  assign T180 = 3'h4 == in_1;
  assign T181 = T187 | T182;
  assign T182 = T236 & T183;
  assign T183 = 3'h2;
  assign T236 = T184 ? 3'h7 : 3'h0;
  assign T184 = T185;
  assign T185 = T186;
  assign T186 = io_config[3'h5];
  assign T187 = T3 & T188;
  assign T188 = ~ T183;
  assign T189 = 3'h5 == in_1;
  assign T190 = T196 | T191;
  assign T191 = T237 & T192;
  assign T192 = 3'h2;
  assign T237 = T193 ? 3'h7 : 3'h0;
  assign T193 = T194;
  assign T194 = T195;
  assign T195 = io_config[3'h6];
  assign T196 = T2 & T197;
  assign T197 = ~ T192;
  assign T198 = 3'h6 == in_1;
  assign T199 = T205 | T200;
  assign T200 = T238 & T201;
  assign T201 = 3'h2;
  assign T238 = T202 ? 3'h7 : 3'h0;
  assign T202 = T203;
  assign T203 = T204;
  assign T204 = io_config[3'h7];
  assign T205 = T1 & T206;
  assign T206 = ~ T201;
  assign T207 = 3'h7 == in_1;
endmodule

module CarryChainModule(
    input [1:0] io_propagate,
    input [1:0] io_generate,
    input  io_carry_in,
    output[1:0] io_out,
    output io_carry_out
);

  wire T0;
  wire T1;
  wire mux0_out;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[1:0] T20;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T21;
  wire T9;
  wire T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T22;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[1:0] T23;
  wire T16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;


  assign io_carry_out = T0;
  assign T0 = T5 ? mux0_out : T1;
  assign T1 = io_generate[1'h1];
  assign mux0_out = T2;
  assign T2 = T4 ? io_carry_in : T3;
  assign T3 = io_generate[1'h0];
  assign T4 = io_propagate[1'h0];
  assign T5 = io_propagate[1'h1];
  assign io_out = T20;
  assign T20 = T6[1'h1:1'h0];
  assign T6 = T11 | T7;
  assign T7 = T21 & T8;
  assign T8 = 3'h2;
  assign T21 = T9 ? 3'h7 : 3'h0;
  assign T9 = T10;
  assign T10 = mux0_out;
  assign T11 = T22 & T12;
  assign T12 = ~ T8;
  assign T22 = {1'h0, T13};
  assign T13 = T18 | T14;
  assign T14 = T23 & T15;
  assign T15 = 2'h1;
  assign T23 = T16 ? 2'h3 : 2'h0;
  assign T16 = T17;
  assign T17 = io_carry_in;
  assign T18 = 2'h0 & T19;
  assign T19 = ~ T15;
endmodule

module ResultFunctionModule(
    input [1:0] io_U,
    input [1:0] io_V,
    input [1:0] io_K,
    input [1:0] io_mx,
    input  io_carry_out,
    output[1:0] io_out
);

  wire[1:0] T26;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T27;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire[1:0] T28;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T29;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T30;
  wire T20;
  wire[2:0] T31;
  wire[1:0] T21;
  wire T22;
  wire[2:0] T32;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;


  assign io_out = T26;
  assign T26 = T0[1'h1:1'h0];
  assign T0 = T25 ? T32 : T1;
  assign T1 = T22 ? T31 : T2;
  assign T2 = T20 ? T13 : T27;
  assign T27 = {1'h0, T3};
  assign T3 = T20 ? T6 : T4;
  assign T4 = T5 ? io_V : 2'h0;
  assign T5 = 2'h0 == io_mx;
  assign T6 = T11 | T7;
  assign T7 = T28 & T8;
  assign T8 = 2'h1;
  assign T28 = T9 ? 2'h3 : 2'h0;
  assign T9 = T10;
  assign T10 = io_carry_out;
  assign T11 = T4 & T12;
  assign T12 = ~ T8;
  assign T13 = T18 | T14;
  assign T14 = T29 & T15;
  assign T15 = 3'h2;
  assign T29 = T16 ? 3'h7 : 3'h0;
  assign T16 = T17;
  assign T17 = io_carry_out;
  assign T18 = T30 & T19;
  assign T19 = ~ T15;
  assign T30 = {1'h0, T3};
  assign T20 = 2'h1 == io_mx;
  assign T31 = {1'h0, T21};
  assign T21 = io_U ^ io_K;
  assign T22 = 2'h2 == io_mx;
  assign T32 = {1'h0, T23};
  assign T23 = ~ T24;
  assign T24 = io_U ^ io_K;
  assign T25 = 2'h3 == io_mx;
endmodule

module TableSelectorModule(
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    input [1:0] io_sel,
    output[1:0] io_out
);

  wire[1:0] T22;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T23;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T24;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T25;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire[1:0] T21;


  assign io_out = T22;
  assign T22 = T0[1'h1:1'h0];
  assign T0 = T9 | T1;
  assign T1 = T23 & T2;
  assign T2 = 3'h2;
  assign T23 = T3 ? 3'h7 : 3'h0;
  assign T3 = T4;
  assign T4 = T5;
  assign T5 = T8 ? T7 : T6;
  assign T6 = io_in_0[1'h1];
  assign T7 = io_in_1[1'h1];
  assign T8 = io_sel[1'h1];
  assign T9 = T24 & T10;
  assign T10 = ~ T2;
  assign T24 = {1'h0, T11};
  assign T11 = T20 | T12;
  assign T12 = T25 & T13;
  assign T13 = 2'h1;
  assign T25 = T14 ? 2'h3 : 2'h0;
  assign T14 = T15;
  assign T15 = T16;
  assign T16 = T19 ? T18 : T17;
  assign T17 = io_in_0[1'h0];
  assign T18 = io_in_1[1'h0];
  assign T19 = io_sel[1'h0];
  assign T20 = 2'h0 & T21;
  assign T21 = ~ T13;
endmodule

module SelectorModule(
    input [1:0] io_in_3,
    input [1:0] io_in_2,
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    input [1:0] io_sel,
    output[1:0] io_out
);

  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_out = T0;
  assign T0 = T7 ? io_in_3 : T1;
  assign T1 = T6 ? io_in_2 : T2;
  assign T2 = T5 ? io_in_1 : T3;
  assign T3 = T4 ? io_in_0 : 2'h2;
  assign T4 = 2'h0 == io_sel;
  assign T5 = 2'h1 == io_sel;
  assign T6 = 2'h2 == io_sel;
  assign T7 = 2'h3 == io_sel;
endmodule

module FunctionalUnitModule(
    input [1:0] io_X_in_3,
    input [1:0] io_X_in_2,
    input [1:0] io_X_in_1,
    input [1:0] io_X_in_0,
    input  io_shift_X_in_2,
    input  io_shift_X_in_1,
    input  io_shift_X_in_0,
    input [1:0] io_H_out_above,
    input  io_shift_carry_in,
    input  io_carry_in,
    input [63:0] io_config,
    output io_shift_X_out_2,
    output io_shift_X_out_1,
    output io_shift_X_out_0,
    output io_shift_carry_out,
    output io_carry_out,
    output[1:0] io_Z
);

  wire[1:0] shiftinvert_out_2;
  wire[1:0] shiftinvert_out_0;
  wire[1:0] shiftinvert_out_1;
  wire[1:0] T0;
  wire T1;
  wire T2;
  wire[1:0] mx;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  wire[1:0] D_sel_out;
  wire[1:0] T7;
  wire[1:0] crossbar_out_3;
  wire D_sel;
  wire T8;
  wire[2:0] mode;
  wire[2:0] T9;
  wire[1:0] lut_out_0;
  wire[1:0] lut_out_1;
  wire[1:0] carrychain_out;
  wire T10;
  wire T11;
  wire T12;
  wire[7:0] T13;
  wire[1:0] lut_in_0;
  wire[1:0] T14;
  wire[1:0] crossbar_out_0;
  wire[1:0] csa_out_carry;
  wire csa_or_crossbar;
  wire T15;
  wire[1:0] T16;
  wire[1:0] lut_in_1;
  wire[1:0] T17;
  wire[1:0] crossbar_out_1;
  wire[1:0] csa_out_sum;
  wire[1:0] lut_in_2;
  wire[1:0] crossbar_out_2;
  wire[7:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire[1:0] X_in_sel_2;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire[1:0] X_in_sel_1;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire[1:0] X_in_sel_0;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire[1:0] X_in_sel_3;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] tableselector_out;
  wire T39;
  wire[1:0] T40;
  wire[1:0] selector_out;
  wire T41;
  wire T42;
  wire[1:0] resultfunct_out;
  wire T43;
  wire[1:0] CrossbarModule_io_out;
  wire[1:0] CrossbarModule_1_io_out;
  wire[1:0] CrossbarModule_2_io_out;
  wire[1:0] CrossbarModule_3_io_out;
  wire[1:0] ShiftInvertModule_io_out;
  wire ShiftInvertModule_io_shift_out;
  wire[1:0] ShiftInvertModule_1_io_out;
  wire ShiftInvertModule_1_io_shift_out;
  wire[1:0] ShiftInvertModule_2_io_out;
  wire ShiftInvertModule_2_io_shift_out;
  wire[1:0] CarrySaveAdderModule_io_sum;
  wire[1:0] CarrySaveAdderModule_io_carry;
  wire CarrySaveAdderModule_io_shift_carry_out;
  wire[1:0] LookUpTableModule_io_out;
  wire[1:0] LookUpTableModule_1_io_out;
  wire[1:0] CarryChainModule_io_out;
  wire CarryChainModule_io_carry_out;
  wire[1:0] ResultFunctionModule_io_out;
  wire[1:0] TableSelectorModule_io_out;
  wire[1:0] SelectorModule_io_out;


  assign shiftinvert_out_2 = ShiftInvertModule_2_io_out;
  assign shiftinvert_out_0 = ShiftInvertModule_io_out;
  assign shiftinvert_out_1 = ShiftInvertModule_1_io_out;
  assign T0 = T1 ? io_X_in_1 : io_X_in_3;
  assign T1 = T2;
  assign T2 = mx[1'h0];
  assign mx = T3;
  assign T3 = io_config[6'h21:6'h20];
  assign T4 = T5 ? 2'h0 : io_H_out_above;
  assign T5 = T6;
  assign T6 = mx[1'h0];
  assign D_sel_out = T7;
  assign T7 = D_sel ? 2'h2 : crossbar_out_3;
  assign crossbar_out_3 = CrossbarModule_3_io_out;
  assign D_sel = T8;
  assign T8 = mode[1'h0];
  assign mode = T9;
  assign T9 = io_config[4'hf:4'hd];
  assign lut_out_0 = LookUpTableModule_io_out;
  assign lut_out_1 = LookUpTableModule_1_io_out;
  assign carrychain_out = CarryChainModule_io_out;
  assign T10 = T11 ? io_carry_in : 1'h0;
  assign T11 = T12;
  assign T12 = mode[1'h0];
  assign T13 = io_config[5'h1f:5'h18];
  assign lut_in_0 = T14;
  assign T14 = csa_or_crossbar ? csa_out_carry : crossbar_out_0;
  assign crossbar_out_0 = CrossbarModule_io_out;
  assign csa_out_carry = CarrySaveAdderModule_io_carry;
  assign csa_or_crossbar = T15;
  assign T15 = T16 == 2'h3;
  assign T16 = mode[2'h2:1'h1];
  assign lut_in_1 = T17;
  assign T17 = csa_or_crossbar ? csa_out_sum : crossbar_out_1;
  assign crossbar_out_1 = CrossbarModule_1_io_out;
  assign csa_out_sum = CarrySaveAdderModule_io_sum;
  assign lut_in_2 = crossbar_out_2;
  assign crossbar_out_2 = CrossbarModule_2_io_out;
  assign T18 = io_config[5'h17:5'h10];
  assign T19 = T20 ? io_shift_carry_in : 1'h0;
  assign T20 = T21;
  assign T21 = mode[1'h0];
  assign X_in_sel_2 = T22;
  assign T22 = io_config[6'h29:6'h28];
  assign T23 = T24 ? io_shift_X_in_2 : 1'h0;
  assign T24 = T25;
  assign T25 = mode[1'h0];
  assign X_in_sel_1 = T26;
  assign T26 = io_config[6'h31:6'h30];
  assign T27 = T28 ? io_shift_X_in_1 : 1'h0;
  assign T28 = T29;
  assign T29 = mode[1'h0];
  assign X_in_sel_0 = T30;
  assign T30 = io_config[6'h39:6'h38];
  assign T31 = T32 ? io_shift_X_in_0 : 1'h0;
  assign T32 = T33;
  assign T33 = mode[1'h0];
  assign X_in_sel_3 = T34;
  assign T34 = io_config[6'h21:6'h20];
  assign io_Z = T35;
  assign T35 = T43 ? resultfunct_out : T36;
  assign T36 = T42 ? resultfunct_out : T37;
  assign T37 = T41 ? selector_out : T38;
  assign T38 = T39 ? tableselector_out : 2'h0;
  assign tableselector_out = TableSelectorModule_io_out;
  assign T39 = 2'h0 == T40;
  assign T40 = mode[2'h2:1'h1];
  assign selector_out = SelectorModule_io_out;
  assign T41 = 2'h1 == T40;
  assign T42 = 2'h2 == T40;
  assign resultfunct_out = ResultFunctionModule_io_out;
  assign T43 = 2'h3 == T40;
  assign io_carry_out = CarryChainModule_io_carry_out;
  assign io_shift_carry_out = CarrySaveAdderModule_io_shift_carry_out;
  assign io_shift_X_out_0 = ShiftInvertModule_io_shift_out;
  assign io_shift_X_out_1 = ShiftInvertModule_1_io_shift_out;
  assign io_shift_X_out_2 = ShiftInvertModule_2_io_shift_out;
  CrossbarModule CrossbarModule(
       .io_in( io_X_in_0 ),
       .io_sel( X_in_sel_0 ),
       .io_out( CrossbarModule_io_out )
  );
  CrossbarModule CrossbarModule_1(
       .io_in( io_X_in_1 ),
       .io_sel( X_in_sel_1 ),
       .io_out( CrossbarModule_1_io_out )
  );
  CrossbarModule CrossbarModule_2(
       .io_in( io_X_in_2 ),
       .io_sel( X_in_sel_2 ),
       .io_out( CrossbarModule_2_io_out )
  );
  CrossbarModule CrossbarModule_3(
       .io_in( io_X_in_3 ),
       .io_sel( X_in_sel_3 ),
       .io_out( CrossbarModule_3_io_out )
  );
  ShiftInvertModule ShiftInvertModule(
       .io_shift_in( T31 ),
       .io_in( io_X_in_0 ),
       .io_sel( X_in_sel_0 ),
       .io_out( ShiftInvertModule_io_out ),
       .io_shift_out( ShiftInvertModule_io_shift_out )
  );
  ShiftInvertModule ShiftInvertModule_1(
       .io_shift_in( T27 ),
       .io_in( io_X_in_1 ),
       .io_sel( X_in_sel_1 ),
       .io_out( ShiftInvertModule_1_io_out ),
       .io_shift_out( ShiftInvertModule_1_io_shift_out )
  );
  ShiftInvertModule ShiftInvertModule_2(
       .io_shift_in( T23 ),
       .io_in( io_X_in_2 ),
       .io_sel( X_in_sel_2 ),
       .io_out( ShiftInvertModule_2_io_out ),
       .io_shift_out( ShiftInvertModule_2_io_shift_out )
  );
  CarrySaveAdderModule CarrySaveAdderModule(
       .io_shift_carry_in( T19 ),
       .io_in_2( shiftinvert_out_2 ),
       .io_in_1( shiftinvert_out_1 ),
       .io_in_0( shiftinvert_out_0 ),
       .io_sum( CarrySaveAdderModule_io_sum ),
       .io_carry( CarrySaveAdderModule_io_carry ),
       .io_shift_carry_out( CarrySaveAdderModule_io_shift_carry_out )
  );
  LookUpTableModule LookUpTableModule(
       .io_in_2( lut_in_2 ),
       .io_in_1( lut_in_1 ),
       .io_in_0( lut_in_0 ),
       .io_config( T18 ),
       .io_out( LookUpTableModule_io_out )
  );
  LookUpTableModule LookUpTableModule_1(
       .io_in_2( lut_in_2 ),
       .io_in_1( lut_in_1 ),
       .io_in_0( lut_in_0 ),
       .io_config( T13 ),
       .io_out( LookUpTableModule_1_io_out )
  );
  CarryChainModule CarryChainModule(
       .io_propagate( lut_out_1 ),
       .io_generate( lut_out_0 ),
       .io_carry_in( T10 ),
       .io_out( CarryChainModule_io_out ),
       .io_carry_out( CarryChainModule_io_carry_out )
  );
  ResultFunctionModule ResultFunctionModule(
       .io_U( lut_out_1 ),
       .io_V( lut_out_0 ),
       .io_K( carrychain_out ),
       .io_mx( mx ),
       .io_carry_out( CarryChainModule_io_carry_out ),
       .io_out( ResultFunctionModule_io_out )
  );
  TableSelectorModule TableSelectorModule(
       .io_in_1( lut_out_1 ),
       .io_in_0( lut_out_0 ),
       .io_sel( D_sel_out ),
       .io_out( TableSelectorModule_io_out )
  );
  SelectorModule SelectorModule(
       .io_in_3( T4 ),
       .io_in_2( T0 ),
       .io_in_1( shiftinvert_out_1 ),
       .io_in_0( shiftinvert_out_0 ),
       .io_sel( shiftinvert_out_2 ),
       .io_out( SelectorModule_io_out )
  );
endmodule

module LogicBlockModule(input clk, input reset,
    input [1:0] io_V_wire_in_15,
    input [1:0] io_V_wire_in_14,
    input [1:0] io_V_wire_in_13,
    input [1:0] io_V_wire_in_12,
    input [1:0] io_V_wire_in_11,
    input [1:0] io_V_wire_in_10,
    input [1:0] io_V_wire_in_9,
    input [1:0] io_V_wire_in_8,
    input [1:0] io_V_wire_in_7,
    input [1:0] io_V_wire_in_6,
    input [1:0] io_V_wire_in_5,
    input [1:0] io_V_wire_in_4,
    input [1:0] io_V_wire_in_3,
    input [1:0] io_V_wire_in_2,
    input [1:0] io_V_wire_in_1,
    input [1:0] io_V_wire_in_0,
    input [1:0] io_H_wire_above_in_10,
    input [1:0] io_H_wire_above_in_9,
    input [1:0] io_H_wire_above_in_8,
    input [1:0] io_H_wire_above_in_7,
    input [1:0] io_H_wire_above_in_6,
    input [1:0] io_H_wire_above_in_5,
    input [1:0] io_H_wire_above_in_4,
    input [1:0] io_H_wire_above_in_3,
    input [1:0] io_H_wire_above_in_2,
    input [1:0] io_H_wire_above_in_1,
    input [1:0] io_H_wire_above_in_0,
    input [1:0] io_H_wire_below_in_10,
    input [1:0] io_H_wire_below_in_9,
    input [1:0] io_H_wire_below_in_8,
    input [1:0] io_H_wire_below_in_7,
    input [1:0] io_H_wire_below_in_6,
    input [1:0] io_H_wire_below_in_5,
    input [1:0] io_H_wire_below_in_4,
    input [1:0] io_H_wire_below_in_3,
    input [1:0] io_H_wire_below_in_2,
    input [1:0] io_H_wire_below_in_1,
    input [1:0] io_H_wire_below_in_0,
    input [1:0] io_G_wire_above_in_3,
    input [1:0] io_G_wire_above_in_2,
    input [1:0] io_G_wire_above_in_1,
    input [1:0] io_G_wire_above_in_0,
    input [1:0] io_G_wire_below_in_3,
    input [1:0] io_G_wire_below_in_2,
    input [1:0] io_G_wire_below_in_1,
    input [1:0] io_G_wire_below_in_0,
    input [1:0] io_mem_bus_in,
    input  io_shift_X_in_2,
    input  io_shift_X_in_1,
    input  io_shift_X_in_0,
    input [1:0] io_H_out_above,
    input  io_shift_carry_in,
    input  io_carry_in,
    output io_shift_X_out_2,
    output io_shift_X_out_1,
    output io_shift_X_out_0,
    output io_shift_carry_out,
    output io_carry_out,
    input  io_store_en,
    input  io_mem_D_or_Z,
    input [63:0] io_config,
    output[1:0] io_mem_bus_out,
    output[1:0] io_V_wire_out,
    output[1:0] io_H_wire_out,
    output[1:0] io_G_wire_out,
    output[2:0] io_config_G_out,
    output[4:0] io_config_V_out
);

  wire[1:0] X_in_0;
  wire[1:0] X_in_1;
  wire[1:0] X_in_2;
  wire[1:0] X_in_3;
  reg [1:0] D_reg;
  wire[1:0] T36;
  wire[1:0] T0;
  wire[1:0] D_reg_in;
  wire[1:0] T1;
  wire T2;
  wire store_D;
  wire T3;
  wire T4;
  wire T5;
  wire D_sel;
  wire T6;
  wire T7;
  reg [1:0] Z_reg;
  wire[1:0] T37;
  wire[1:0] T8;
  wire[1:0] Z_reg_in;
  wire[1:0] T9;
  wire[1:0] Z;
  wire T10;
  wire store_Z;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire Z_sel;
  wire T15;
  wire T16;
  wire[5:0] config_X_in_0;
  wire[5:0] T17;
  wire[5:0] config_X_in_1;
  wire[5:0] T18;
  wire[5:0] config_X_in_2;
  wire[5:0] T19;
  wire[5:0] config_X_in_3;
  wire[5:0] T20;
  wire[4:0] T21;
  wire[2:0] T22;
  wire[1:0] T23;
  wire[1:0] Z_out;
  wire[1:0] T24;
  wire[1:0] D_out;
  wire[1:0] T25;
  wire G_sel;
  wire T26;
  wire T27;
  wire[1:0] T28;
  wire H_sel;
  wire T29;
  wire T30;
  wire[1:0] T31;
  wire V_sel;
  wire T32;
  wire T33;
  wire[1:0] T34;
  wire T35;
  wire[1:0] LogicBlockInBBModule_io_X_in_3;
  wire[1:0] LogicBlockInBBModule_io_X_in_2;
  wire[1:0] LogicBlockInBBModule_io_X_in_1;
  wire[1:0] LogicBlockInBBModule_io_X_in_0;
  wire FUpeek_io_shift_X_out_2;
  wire FUpeek_io_shift_X_out_1;
  wire FUpeek_io_shift_X_out_0;
  wire FUpeek_io_shift_carry_out;
  wire FUpeek_io_carry_out;
  wire[1:0] FUpeek_io_Z;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    D_reg = {1{$random}};
    Z_reg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign X_in_0 = LogicBlockInBBModule_io_X_in_0;
  assign X_in_1 = LogicBlockInBBModule_io_X_in_1;
  assign X_in_2 = LogicBlockInBBModule_io_X_in_2;
  assign X_in_3 = LogicBlockInBBModule_io_X_in_3;
  assign T36 = reset ? 2'h0 : T0;
  assign T0 = T4 ? D_reg_in : D_reg;
  assign D_reg_in = T1;
  assign T1 = T2 ? io_mem_bus_in : X_in_3;
  assign T2 = store_D;
  assign store_D = T3;
  assign T3 = io_store_en & io_mem_D_or_Z;
  assign T4 = D_sel | T5;
  assign T5 = store_D;
  assign D_sel = T6;
  assign T6 = T7;
  assign T7 = io_config[4'hb];
  assign T37 = reset ? 2'h0 : T8;
  assign T8 = T13 ? Z_reg_in : Z_reg;
  assign Z_reg_in = T9;
  assign T9 = T10 ? io_mem_bus_in : Z;
  assign Z = FUpeek_io_Z;
  assign T10 = store_Z;
  assign store_Z = T11;
  assign T11 = io_store_en & T12;
  assign T12 = ~ io_mem_D_or_Z;
  assign T13 = Z_sel | T14;
  assign T14 = store_Z;
  assign Z_sel = T15;
  assign T15 = T16;
  assign T16 = io_config[4'hc];
  assign config_X_in_0 = T17;
  assign T17 = io_config[6'h3f:6'h3a];
  assign config_X_in_1 = T18;
  assign T18 = io_config[6'h37:6'h32];
  assign config_X_in_2 = T19;
  assign T19 = io_config[6'h2f:6'h2a];
  assign config_X_in_3 = T20;
  assign T20 = io_config[6'h27:6'h22];
  assign io_config_V_out = T21;
  assign T21 = io_config[3'h4:1'h0];
  assign io_config_G_out = T22;
  assign T22 = io_config[3'h7:3'h5];
  assign io_G_wire_out = T23;
  assign T23 = G_sel ? D_out : Z_out;
  assign Z_out = T24;
  assign T24 = Z_sel ? Z_reg : Z;
  assign D_out = T25;
  assign T25 = D_sel ? D_reg : X_in_3;
  assign G_sel = T26;
  assign T26 = T27;
  assign T27 = io_config[4'h9];
  assign io_H_wire_out = T28;
  assign T28 = H_sel ? D_out : Z_out;
  assign H_sel = T29;
  assign T29 = T30;
  assign T30 = io_config[4'ha];
  assign io_V_wire_out = T31;
  assign T31 = V_sel ? D_out : Z_out;
  assign V_sel = T32;
  assign T32 = T33;
  assign T33 = io_config[4'h8];
  assign io_mem_bus_out = T34;
  assign T34 = T35 ? D_reg : Z_reg;
  assign T35 = io_mem_D_or_Z;
  assign io_carry_out = FUpeek_io_carry_out;
  assign io_shift_carry_out = FUpeek_io_shift_carry_out;
  assign io_shift_X_out_0 = FUpeek_io_shift_X_out_0;
  assign io_shift_X_out_1 = FUpeek_io_shift_X_out_1;
  assign io_shift_X_out_2 = FUpeek_io_shift_X_out_2;
  LogicBlockInBBModule LogicBlockInBBModule(
       .io_V_wire_in_15( io_V_wire_in_15 ),
       .io_V_wire_in_14( io_V_wire_in_14 ),
       .io_V_wire_in_13( io_V_wire_in_13 ),
       .io_V_wire_in_12( io_V_wire_in_12 ),
       .io_V_wire_in_11( io_V_wire_in_11 ),
       .io_V_wire_in_10( io_V_wire_in_10 ),
       .io_V_wire_in_9( io_V_wire_in_9 ),
       .io_V_wire_in_8( io_V_wire_in_8 ),
       .io_V_wire_in_7( io_V_wire_in_7 ),
       .io_V_wire_in_6( io_V_wire_in_6 ),
       .io_V_wire_in_5( io_V_wire_in_5 ),
       .io_V_wire_in_4( io_V_wire_in_4 ),
       .io_V_wire_in_3( io_V_wire_in_3 ),
       .io_V_wire_in_2( io_V_wire_in_2 ),
       .io_V_wire_in_1( io_V_wire_in_1 ),
       .io_V_wire_in_0( io_V_wire_in_0 ),
       .io_H_wire_above_in_10( io_H_wire_above_in_10 ),
       .io_H_wire_above_in_9( io_H_wire_above_in_9 ),
       .io_H_wire_above_in_8( io_H_wire_above_in_8 ),
       .io_H_wire_above_in_7( io_H_wire_above_in_7 ),
       .io_H_wire_above_in_6( io_H_wire_above_in_6 ),
       .io_H_wire_above_in_5( io_H_wire_above_in_5 ),
       .io_H_wire_above_in_4( io_H_wire_above_in_4 ),
       .io_H_wire_above_in_3( io_H_wire_above_in_3 ),
       .io_H_wire_above_in_2( io_H_wire_above_in_2 ),
       .io_H_wire_above_in_1( io_H_wire_above_in_1 ),
       .io_H_wire_above_in_0( io_H_wire_above_in_0 ),
       .io_H_wire_below_in_10( io_H_wire_below_in_10 ),
       .io_H_wire_below_in_9( io_H_wire_below_in_9 ),
       .io_H_wire_below_in_8( io_H_wire_below_in_8 ),
       .io_H_wire_below_in_7( io_H_wire_below_in_7 ),
       .io_H_wire_below_in_6( io_H_wire_below_in_6 ),
       .io_H_wire_below_in_5( io_H_wire_below_in_5 ),
       .io_H_wire_below_in_4( io_H_wire_below_in_4 ),
       .io_H_wire_below_in_3( io_H_wire_below_in_3 ),
       .io_H_wire_below_in_2( io_H_wire_below_in_2 ),
       .io_H_wire_below_in_1( io_H_wire_below_in_1 ),
       .io_H_wire_below_in_0( io_H_wire_below_in_0 ),
       .io_G_wire_above_in_3( io_G_wire_above_in_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_in_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_in_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_in_0 ),
       .io_G_wire_below_in_3( io_G_wire_below_in_3 ),
       .io_G_wire_below_in_2( io_G_wire_below_in_2 ),
       .io_G_wire_below_in_1( io_G_wire_below_in_1 ),
       .io_G_wire_below_in_0( io_G_wire_below_in_0 ),
       .io_config_X_in_3( config_X_in_3 ),
       .io_config_X_in_2( config_X_in_2 ),
       .io_config_X_in_1( config_X_in_1 ),
       .io_config_X_in_0( config_X_in_0 ),
       .io_Z_reg( Z_reg ),
       .io_D_reg( D_reg ),
       .io_X_in_3( LogicBlockInBBModule_io_X_in_3 ),
       .io_X_in_2( LogicBlockInBBModule_io_X_in_2 ),
       .io_X_in_1( LogicBlockInBBModule_io_X_in_1 ),
       .io_X_in_0( LogicBlockInBBModule_io_X_in_0 )
  );
  FunctionalUnitModule FUpeek(
       .io_X_in_3( X_in_3 ),
       .io_X_in_2( X_in_2 ),
       .io_X_in_1( X_in_1 ),
       .io_X_in_0( X_in_0 ),
       .io_shift_X_in_2( io_shift_X_in_2 ),
       .io_shift_X_in_1( io_shift_X_in_1 ),
       .io_shift_X_in_0( io_shift_X_in_0 ),
       .io_H_out_above( io_H_out_above ),
       .io_shift_carry_in( io_shift_carry_in ),
       .io_carry_in( io_carry_in ),
       .io_config( io_config ),
       .io_shift_X_out_2( FUpeek_io_shift_X_out_2 ),
       .io_shift_X_out_1( FUpeek_io_shift_X_out_1 ),
       .io_shift_X_out_0( FUpeek_io_shift_X_out_0 ),
       .io_shift_carry_out( FUpeek_io_shift_carry_out ),
       .io_carry_out( FUpeek_io_carry_out ),
       .io_Z( FUpeek_io_Z )
  );

  always @(posedge clk) begin
    if(reset) begin
      D_reg <= 2'h0;
    end else if(T4) begin
      D_reg <= D_reg_in;
    end
    if(reset) begin
      Z_reg <= 2'h0;
    end else if(T13) begin
      Z_reg <= Z_reg_in;
    end
  end
endmodule

module GWireModule(
    input [1:0] io_G_in_22,
    input [1:0] io_G_in_21,
    input [1:0] io_G_in_20,
    input [1:0] io_G_in_19,
    input [1:0] io_G_in_18,
    input [1:0] io_G_in_17,
    input [1:0] io_G_in_16,
    input [1:0] io_G_in_15,
    input [1:0] io_G_in_14,
    input [1:0] io_G_in_13,
    input [1:0] io_G_in_12,
    input [1:0] io_G_in_11,
    input [1:0] io_G_in_10,
    input [1:0] io_G_in_9,
    input [1:0] io_G_in_8,
    input [1:0] io_G_in_7,
    input [1:0] io_G_in_6,
    input [1:0] io_G_in_5,
    input [1:0] io_G_in_4,
    input [1:0] io_G_in_3,
    input [1:0] io_G_in_2,
    input [1:0] io_G_in_1,
    input [1:0] io_G_in_0,
    input [22:0] io_en,
    output[1:0] io_G_out
);

  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;


  assign io_G_out = T0;
  assign T0 = T67 ? io_G_in_22 : T1;
  assign T1 = T65 ? io_G_in_21 : T2;
  assign T2 = T63 ? io_G_in_20 : T3;
  assign T3 = T61 ? io_G_in_19 : T4;
  assign T4 = T59 ? io_G_in_18 : T5;
  assign T5 = T57 ? io_G_in_17 : T6;
  assign T6 = T55 ? io_G_in_16 : T7;
  assign T7 = T53 ? io_G_in_15 : T8;
  assign T8 = T51 ? io_G_in_14 : T9;
  assign T9 = T49 ? io_G_in_13 : T10;
  assign T10 = T47 ? io_G_in_12 : T11;
  assign T11 = T45 ? io_G_in_11 : T12;
  assign T12 = T43 ? io_G_in_10 : T13;
  assign T13 = T41 ? io_G_in_9 : T14;
  assign T14 = T39 ? io_G_in_8 : T15;
  assign T15 = T37 ? io_G_in_7 : T16;
  assign T16 = T35 ? io_G_in_6 : T17;
  assign T17 = T33 ? io_G_in_5 : T18;
  assign T18 = T31 ? io_G_in_4 : T19;
  assign T19 = T29 ? io_G_in_3 : T20;
  assign T20 = T27 ? io_G_in_2 : T21;
  assign T21 = T25 ? io_G_in_1 : T22;
  assign T22 = T23 ? io_G_in_0 : 2'h0;
  assign T23 = T24;
  assign T24 = io_en[1'h0];
  assign T25 = T26;
  assign T26 = io_en[1'h1];
  assign T27 = T28;
  assign T28 = io_en[2'h2];
  assign T29 = T30;
  assign T30 = io_en[2'h3];
  assign T31 = T32;
  assign T32 = io_en[3'h4];
  assign T33 = T34;
  assign T34 = io_en[3'h5];
  assign T35 = T36;
  assign T36 = io_en[3'h6];
  assign T37 = T38;
  assign T38 = io_en[3'h7];
  assign T39 = T40;
  assign T40 = io_en[4'h8];
  assign T41 = T42;
  assign T42 = io_en[4'h9];
  assign T43 = T44;
  assign T44 = io_en[4'ha];
  assign T45 = T46;
  assign T46 = io_en[4'hb];
  assign T47 = T48;
  assign T48 = io_en[4'hc];
  assign T49 = T50;
  assign T50 = io_en[4'hd];
  assign T51 = T52;
  assign T52 = io_en[4'he];
  assign T53 = T54;
  assign T54 = io_en[4'hf];
  assign T55 = T56;
  assign T56 = io_en[5'h10];
  assign T57 = T58;
  assign T58 = io_en[5'h11];
  assign T59 = T60;
  assign T60 = io_en[5'h12];
  assign T61 = T62;
  assign T62 = io_en[5'h13];
  assign T63 = T64;
  assign T64 = io_en[5'h14];
  assign T65 = T66;
  assign T66 = io_en[5'h15];
  assign T67 = T68;
  assign T68 = io_en[5'h16];
endmodule

module ArrayRowModule(input clk, input reset,
    input [1:0] io_V_wire_in_367,
    input [1:0] io_V_wire_in_366,
    input [1:0] io_V_wire_in_365,
    input [1:0] io_V_wire_in_364,
    input [1:0] io_V_wire_in_363,
    input [1:0] io_V_wire_in_362,
    input [1:0] io_V_wire_in_361,
    input [1:0] io_V_wire_in_360,
    input [1:0] io_V_wire_in_359,
    input [1:0] io_V_wire_in_358,
    input [1:0] io_V_wire_in_357,
    input [1:0] io_V_wire_in_356,
    input [1:0] io_V_wire_in_355,
    input [1:0] io_V_wire_in_354,
    input [1:0] io_V_wire_in_353,
    input [1:0] io_V_wire_in_352,
    input [1:0] io_V_wire_in_351,
    input [1:0] io_V_wire_in_350,
    input [1:0] io_V_wire_in_349,
    input [1:0] io_V_wire_in_348,
    input [1:0] io_V_wire_in_347,
    input [1:0] io_V_wire_in_346,
    input [1:0] io_V_wire_in_345,
    input [1:0] io_V_wire_in_344,
    input [1:0] io_V_wire_in_343,
    input [1:0] io_V_wire_in_342,
    input [1:0] io_V_wire_in_341,
    input [1:0] io_V_wire_in_340,
    input [1:0] io_V_wire_in_339,
    input [1:0] io_V_wire_in_338,
    input [1:0] io_V_wire_in_337,
    input [1:0] io_V_wire_in_336,
    input [1:0] io_V_wire_in_335,
    input [1:0] io_V_wire_in_334,
    input [1:0] io_V_wire_in_333,
    input [1:0] io_V_wire_in_332,
    input [1:0] io_V_wire_in_331,
    input [1:0] io_V_wire_in_330,
    input [1:0] io_V_wire_in_329,
    input [1:0] io_V_wire_in_328,
    input [1:0] io_V_wire_in_327,
    input [1:0] io_V_wire_in_326,
    input [1:0] io_V_wire_in_325,
    input [1:0] io_V_wire_in_324,
    input [1:0] io_V_wire_in_323,
    input [1:0] io_V_wire_in_322,
    input [1:0] io_V_wire_in_321,
    input [1:0] io_V_wire_in_320,
    input [1:0] io_V_wire_in_319,
    input [1:0] io_V_wire_in_318,
    input [1:0] io_V_wire_in_317,
    input [1:0] io_V_wire_in_316,
    input [1:0] io_V_wire_in_315,
    input [1:0] io_V_wire_in_314,
    input [1:0] io_V_wire_in_313,
    input [1:0] io_V_wire_in_312,
    input [1:0] io_V_wire_in_311,
    input [1:0] io_V_wire_in_310,
    input [1:0] io_V_wire_in_309,
    input [1:0] io_V_wire_in_308,
    input [1:0] io_V_wire_in_307,
    input [1:0] io_V_wire_in_306,
    input [1:0] io_V_wire_in_305,
    input [1:0] io_V_wire_in_304,
    input [1:0] io_V_wire_in_303,
    input [1:0] io_V_wire_in_302,
    input [1:0] io_V_wire_in_301,
    input [1:0] io_V_wire_in_300,
    input [1:0] io_V_wire_in_299,
    input [1:0] io_V_wire_in_298,
    input [1:0] io_V_wire_in_297,
    input [1:0] io_V_wire_in_296,
    input [1:0] io_V_wire_in_295,
    input [1:0] io_V_wire_in_294,
    input [1:0] io_V_wire_in_293,
    input [1:0] io_V_wire_in_292,
    input [1:0] io_V_wire_in_291,
    input [1:0] io_V_wire_in_290,
    input [1:0] io_V_wire_in_289,
    input [1:0] io_V_wire_in_288,
    input [1:0] io_V_wire_in_287,
    input [1:0] io_V_wire_in_286,
    input [1:0] io_V_wire_in_285,
    input [1:0] io_V_wire_in_284,
    input [1:0] io_V_wire_in_283,
    input [1:0] io_V_wire_in_282,
    input [1:0] io_V_wire_in_281,
    input [1:0] io_V_wire_in_280,
    input [1:0] io_V_wire_in_279,
    input [1:0] io_V_wire_in_278,
    input [1:0] io_V_wire_in_277,
    input [1:0] io_V_wire_in_276,
    input [1:0] io_V_wire_in_275,
    input [1:0] io_V_wire_in_274,
    input [1:0] io_V_wire_in_273,
    input [1:0] io_V_wire_in_272,
    input [1:0] io_V_wire_in_271,
    input [1:0] io_V_wire_in_270,
    input [1:0] io_V_wire_in_269,
    input [1:0] io_V_wire_in_268,
    input [1:0] io_V_wire_in_267,
    input [1:0] io_V_wire_in_266,
    input [1:0] io_V_wire_in_265,
    input [1:0] io_V_wire_in_264,
    input [1:0] io_V_wire_in_263,
    input [1:0] io_V_wire_in_262,
    input [1:0] io_V_wire_in_261,
    input [1:0] io_V_wire_in_260,
    input [1:0] io_V_wire_in_259,
    input [1:0] io_V_wire_in_258,
    input [1:0] io_V_wire_in_257,
    input [1:0] io_V_wire_in_256,
    input [1:0] io_V_wire_in_255,
    input [1:0] io_V_wire_in_254,
    input [1:0] io_V_wire_in_253,
    input [1:0] io_V_wire_in_252,
    input [1:0] io_V_wire_in_251,
    input [1:0] io_V_wire_in_250,
    input [1:0] io_V_wire_in_249,
    input [1:0] io_V_wire_in_248,
    input [1:0] io_V_wire_in_247,
    input [1:0] io_V_wire_in_246,
    input [1:0] io_V_wire_in_245,
    input [1:0] io_V_wire_in_244,
    input [1:0] io_V_wire_in_243,
    input [1:0] io_V_wire_in_242,
    input [1:0] io_V_wire_in_241,
    input [1:0] io_V_wire_in_240,
    input [1:0] io_V_wire_in_239,
    input [1:0] io_V_wire_in_238,
    input [1:0] io_V_wire_in_237,
    input [1:0] io_V_wire_in_236,
    input [1:0] io_V_wire_in_235,
    input [1:0] io_V_wire_in_234,
    input [1:0] io_V_wire_in_233,
    input [1:0] io_V_wire_in_232,
    input [1:0] io_V_wire_in_231,
    input [1:0] io_V_wire_in_230,
    input [1:0] io_V_wire_in_229,
    input [1:0] io_V_wire_in_228,
    input [1:0] io_V_wire_in_227,
    input [1:0] io_V_wire_in_226,
    input [1:0] io_V_wire_in_225,
    input [1:0] io_V_wire_in_224,
    input [1:0] io_V_wire_in_223,
    input [1:0] io_V_wire_in_222,
    input [1:0] io_V_wire_in_221,
    input [1:0] io_V_wire_in_220,
    input [1:0] io_V_wire_in_219,
    input [1:0] io_V_wire_in_218,
    input [1:0] io_V_wire_in_217,
    input [1:0] io_V_wire_in_216,
    input [1:0] io_V_wire_in_215,
    input [1:0] io_V_wire_in_214,
    input [1:0] io_V_wire_in_213,
    input [1:0] io_V_wire_in_212,
    input [1:0] io_V_wire_in_211,
    input [1:0] io_V_wire_in_210,
    input [1:0] io_V_wire_in_209,
    input [1:0] io_V_wire_in_208,
    input [1:0] io_V_wire_in_207,
    input [1:0] io_V_wire_in_206,
    input [1:0] io_V_wire_in_205,
    input [1:0] io_V_wire_in_204,
    input [1:0] io_V_wire_in_203,
    input [1:0] io_V_wire_in_202,
    input [1:0] io_V_wire_in_201,
    input [1:0] io_V_wire_in_200,
    input [1:0] io_V_wire_in_199,
    input [1:0] io_V_wire_in_198,
    input [1:0] io_V_wire_in_197,
    input [1:0] io_V_wire_in_196,
    input [1:0] io_V_wire_in_195,
    input [1:0] io_V_wire_in_194,
    input [1:0] io_V_wire_in_193,
    input [1:0] io_V_wire_in_192,
    input [1:0] io_V_wire_in_191,
    input [1:0] io_V_wire_in_190,
    input [1:0] io_V_wire_in_189,
    input [1:0] io_V_wire_in_188,
    input [1:0] io_V_wire_in_187,
    input [1:0] io_V_wire_in_186,
    input [1:0] io_V_wire_in_185,
    input [1:0] io_V_wire_in_184,
    input [1:0] io_V_wire_in_183,
    input [1:0] io_V_wire_in_182,
    input [1:0] io_V_wire_in_181,
    input [1:0] io_V_wire_in_180,
    input [1:0] io_V_wire_in_179,
    input [1:0] io_V_wire_in_178,
    input [1:0] io_V_wire_in_177,
    input [1:0] io_V_wire_in_176,
    input [1:0] io_V_wire_in_175,
    input [1:0] io_V_wire_in_174,
    input [1:0] io_V_wire_in_173,
    input [1:0] io_V_wire_in_172,
    input [1:0] io_V_wire_in_171,
    input [1:0] io_V_wire_in_170,
    input [1:0] io_V_wire_in_169,
    input [1:0] io_V_wire_in_168,
    input [1:0] io_V_wire_in_167,
    input [1:0] io_V_wire_in_166,
    input [1:0] io_V_wire_in_165,
    input [1:0] io_V_wire_in_164,
    input [1:0] io_V_wire_in_163,
    input [1:0] io_V_wire_in_162,
    input [1:0] io_V_wire_in_161,
    input [1:0] io_V_wire_in_160,
    input [1:0] io_V_wire_in_159,
    input [1:0] io_V_wire_in_158,
    input [1:0] io_V_wire_in_157,
    input [1:0] io_V_wire_in_156,
    input [1:0] io_V_wire_in_155,
    input [1:0] io_V_wire_in_154,
    input [1:0] io_V_wire_in_153,
    input [1:0] io_V_wire_in_152,
    input [1:0] io_V_wire_in_151,
    input [1:0] io_V_wire_in_150,
    input [1:0] io_V_wire_in_149,
    input [1:0] io_V_wire_in_148,
    input [1:0] io_V_wire_in_147,
    input [1:0] io_V_wire_in_146,
    input [1:0] io_V_wire_in_145,
    input [1:0] io_V_wire_in_144,
    input [1:0] io_V_wire_in_143,
    input [1:0] io_V_wire_in_142,
    input [1:0] io_V_wire_in_141,
    input [1:0] io_V_wire_in_140,
    input [1:0] io_V_wire_in_139,
    input [1:0] io_V_wire_in_138,
    input [1:0] io_V_wire_in_137,
    input [1:0] io_V_wire_in_136,
    input [1:0] io_V_wire_in_135,
    input [1:0] io_V_wire_in_134,
    input [1:0] io_V_wire_in_133,
    input [1:0] io_V_wire_in_132,
    input [1:0] io_V_wire_in_131,
    input [1:0] io_V_wire_in_130,
    input [1:0] io_V_wire_in_129,
    input [1:0] io_V_wire_in_128,
    input [1:0] io_V_wire_in_127,
    input [1:0] io_V_wire_in_126,
    input [1:0] io_V_wire_in_125,
    input [1:0] io_V_wire_in_124,
    input [1:0] io_V_wire_in_123,
    input [1:0] io_V_wire_in_122,
    input [1:0] io_V_wire_in_121,
    input [1:0] io_V_wire_in_120,
    input [1:0] io_V_wire_in_119,
    input [1:0] io_V_wire_in_118,
    input [1:0] io_V_wire_in_117,
    input [1:0] io_V_wire_in_116,
    input [1:0] io_V_wire_in_115,
    input [1:0] io_V_wire_in_114,
    input [1:0] io_V_wire_in_113,
    input [1:0] io_V_wire_in_112,
    input [1:0] io_V_wire_in_111,
    input [1:0] io_V_wire_in_110,
    input [1:0] io_V_wire_in_109,
    input [1:0] io_V_wire_in_108,
    input [1:0] io_V_wire_in_107,
    input [1:0] io_V_wire_in_106,
    input [1:0] io_V_wire_in_105,
    input [1:0] io_V_wire_in_104,
    input [1:0] io_V_wire_in_103,
    input [1:0] io_V_wire_in_102,
    input [1:0] io_V_wire_in_101,
    input [1:0] io_V_wire_in_100,
    input [1:0] io_V_wire_in_99,
    input [1:0] io_V_wire_in_98,
    input [1:0] io_V_wire_in_97,
    input [1:0] io_V_wire_in_96,
    input [1:0] io_V_wire_in_95,
    input [1:0] io_V_wire_in_94,
    input [1:0] io_V_wire_in_93,
    input [1:0] io_V_wire_in_92,
    input [1:0] io_V_wire_in_91,
    input [1:0] io_V_wire_in_90,
    input [1:0] io_V_wire_in_89,
    input [1:0] io_V_wire_in_88,
    input [1:0] io_V_wire_in_87,
    input [1:0] io_V_wire_in_86,
    input [1:0] io_V_wire_in_85,
    input [1:0] io_V_wire_in_84,
    input [1:0] io_V_wire_in_83,
    input [1:0] io_V_wire_in_82,
    input [1:0] io_V_wire_in_81,
    input [1:0] io_V_wire_in_80,
    input [1:0] io_V_wire_in_79,
    input [1:0] io_V_wire_in_78,
    input [1:0] io_V_wire_in_77,
    input [1:0] io_V_wire_in_76,
    input [1:0] io_V_wire_in_75,
    input [1:0] io_V_wire_in_74,
    input [1:0] io_V_wire_in_73,
    input [1:0] io_V_wire_in_72,
    input [1:0] io_V_wire_in_71,
    input [1:0] io_V_wire_in_70,
    input [1:0] io_V_wire_in_69,
    input [1:0] io_V_wire_in_68,
    input [1:0] io_V_wire_in_67,
    input [1:0] io_V_wire_in_66,
    input [1:0] io_V_wire_in_65,
    input [1:0] io_V_wire_in_64,
    input [1:0] io_V_wire_in_63,
    input [1:0] io_V_wire_in_62,
    input [1:0] io_V_wire_in_61,
    input [1:0] io_V_wire_in_60,
    input [1:0] io_V_wire_in_59,
    input [1:0] io_V_wire_in_58,
    input [1:0] io_V_wire_in_57,
    input [1:0] io_V_wire_in_56,
    input [1:0] io_V_wire_in_55,
    input [1:0] io_V_wire_in_54,
    input [1:0] io_V_wire_in_53,
    input [1:0] io_V_wire_in_52,
    input [1:0] io_V_wire_in_51,
    input [1:0] io_V_wire_in_50,
    input [1:0] io_V_wire_in_49,
    input [1:0] io_V_wire_in_48,
    input [1:0] io_V_wire_in_47,
    input [1:0] io_V_wire_in_46,
    input [1:0] io_V_wire_in_45,
    input [1:0] io_V_wire_in_44,
    input [1:0] io_V_wire_in_43,
    input [1:0] io_V_wire_in_42,
    input [1:0] io_V_wire_in_41,
    input [1:0] io_V_wire_in_40,
    input [1:0] io_V_wire_in_39,
    input [1:0] io_V_wire_in_38,
    input [1:0] io_V_wire_in_37,
    input [1:0] io_V_wire_in_36,
    input [1:0] io_V_wire_in_35,
    input [1:0] io_V_wire_in_34,
    input [1:0] io_V_wire_in_33,
    input [1:0] io_V_wire_in_32,
    input [1:0] io_V_wire_in_31,
    input [1:0] io_V_wire_in_30,
    input [1:0] io_V_wire_in_29,
    input [1:0] io_V_wire_in_28,
    input [1:0] io_V_wire_in_27,
    input [1:0] io_V_wire_in_26,
    input [1:0] io_V_wire_in_25,
    input [1:0] io_V_wire_in_24,
    input [1:0] io_V_wire_in_23,
    input [1:0] io_V_wire_in_22,
    input [1:0] io_V_wire_in_21,
    input [1:0] io_V_wire_in_20,
    input [1:0] io_V_wire_in_19,
    input [1:0] io_V_wire_in_18,
    input [1:0] io_V_wire_in_17,
    input [1:0] io_V_wire_in_16,
    input [1:0] io_V_wire_in_15,
    input [1:0] io_V_wire_in_14,
    input [1:0] io_V_wire_in_13,
    input [1:0] io_V_wire_in_12,
    input [1:0] io_V_wire_in_11,
    input [1:0] io_V_wire_in_10,
    input [1:0] io_V_wire_in_9,
    input [1:0] io_V_wire_in_8,
    input [1:0] io_V_wire_in_7,
    input [1:0] io_V_wire_in_6,
    input [1:0] io_V_wire_in_5,
    input [1:0] io_V_wire_in_4,
    input [1:0] io_V_wire_in_3,
    input [1:0] io_V_wire_in_2,
    input [1:0] io_V_wire_in_1,
    input [1:0] io_V_wire_in_0,
    output[1:0] io_V_wire_out_367,
    output[1:0] io_V_wire_out_366,
    output[1:0] io_V_wire_out_365,
    output[1:0] io_V_wire_out_364,
    output[1:0] io_V_wire_out_363,
    output[1:0] io_V_wire_out_362,
    output[1:0] io_V_wire_out_361,
    output[1:0] io_V_wire_out_360,
    output[1:0] io_V_wire_out_359,
    output[1:0] io_V_wire_out_358,
    output[1:0] io_V_wire_out_357,
    output[1:0] io_V_wire_out_356,
    output[1:0] io_V_wire_out_355,
    output[1:0] io_V_wire_out_354,
    output[1:0] io_V_wire_out_353,
    output[1:0] io_V_wire_out_352,
    output[1:0] io_V_wire_out_351,
    output[1:0] io_V_wire_out_350,
    output[1:0] io_V_wire_out_349,
    output[1:0] io_V_wire_out_348,
    output[1:0] io_V_wire_out_347,
    output[1:0] io_V_wire_out_346,
    output[1:0] io_V_wire_out_345,
    output[1:0] io_V_wire_out_344,
    output[1:0] io_V_wire_out_343,
    output[1:0] io_V_wire_out_342,
    output[1:0] io_V_wire_out_341,
    output[1:0] io_V_wire_out_340,
    output[1:0] io_V_wire_out_339,
    output[1:0] io_V_wire_out_338,
    output[1:0] io_V_wire_out_337,
    output[1:0] io_V_wire_out_336,
    output[1:0] io_V_wire_out_335,
    output[1:0] io_V_wire_out_334,
    output[1:0] io_V_wire_out_333,
    output[1:0] io_V_wire_out_332,
    output[1:0] io_V_wire_out_331,
    output[1:0] io_V_wire_out_330,
    output[1:0] io_V_wire_out_329,
    output[1:0] io_V_wire_out_328,
    output[1:0] io_V_wire_out_327,
    output[1:0] io_V_wire_out_326,
    output[1:0] io_V_wire_out_325,
    output[1:0] io_V_wire_out_324,
    output[1:0] io_V_wire_out_323,
    output[1:0] io_V_wire_out_322,
    output[1:0] io_V_wire_out_321,
    output[1:0] io_V_wire_out_320,
    output[1:0] io_V_wire_out_319,
    output[1:0] io_V_wire_out_318,
    output[1:0] io_V_wire_out_317,
    output[1:0] io_V_wire_out_316,
    output[1:0] io_V_wire_out_315,
    output[1:0] io_V_wire_out_314,
    output[1:0] io_V_wire_out_313,
    output[1:0] io_V_wire_out_312,
    output[1:0] io_V_wire_out_311,
    output[1:0] io_V_wire_out_310,
    output[1:0] io_V_wire_out_309,
    output[1:0] io_V_wire_out_308,
    output[1:0] io_V_wire_out_307,
    output[1:0] io_V_wire_out_306,
    output[1:0] io_V_wire_out_305,
    output[1:0] io_V_wire_out_304,
    output[1:0] io_V_wire_out_303,
    output[1:0] io_V_wire_out_302,
    output[1:0] io_V_wire_out_301,
    output[1:0] io_V_wire_out_300,
    output[1:0] io_V_wire_out_299,
    output[1:0] io_V_wire_out_298,
    output[1:0] io_V_wire_out_297,
    output[1:0] io_V_wire_out_296,
    output[1:0] io_V_wire_out_295,
    output[1:0] io_V_wire_out_294,
    output[1:0] io_V_wire_out_293,
    output[1:0] io_V_wire_out_292,
    output[1:0] io_V_wire_out_291,
    output[1:0] io_V_wire_out_290,
    output[1:0] io_V_wire_out_289,
    output[1:0] io_V_wire_out_288,
    output[1:0] io_V_wire_out_287,
    output[1:0] io_V_wire_out_286,
    output[1:0] io_V_wire_out_285,
    output[1:0] io_V_wire_out_284,
    output[1:0] io_V_wire_out_283,
    output[1:0] io_V_wire_out_282,
    output[1:0] io_V_wire_out_281,
    output[1:0] io_V_wire_out_280,
    output[1:0] io_V_wire_out_279,
    output[1:0] io_V_wire_out_278,
    output[1:0] io_V_wire_out_277,
    output[1:0] io_V_wire_out_276,
    output[1:0] io_V_wire_out_275,
    output[1:0] io_V_wire_out_274,
    output[1:0] io_V_wire_out_273,
    output[1:0] io_V_wire_out_272,
    output[1:0] io_V_wire_out_271,
    output[1:0] io_V_wire_out_270,
    output[1:0] io_V_wire_out_269,
    output[1:0] io_V_wire_out_268,
    output[1:0] io_V_wire_out_267,
    output[1:0] io_V_wire_out_266,
    output[1:0] io_V_wire_out_265,
    output[1:0] io_V_wire_out_264,
    output[1:0] io_V_wire_out_263,
    output[1:0] io_V_wire_out_262,
    output[1:0] io_V_wire_out_261,
    output[1:0] io_V_wire_out_260,
    output[1:0] io_V_wire_out_259,
    output[1:0] io_V_wire_out_258,
    output[1:0] io_V_wire_out_257,
    output[1:0] io_V_wire_out_256,
    output[1:0] io_V_wire_out_255,
    output[1:0] io_V_wire_out_254,
    output[1:0] io_V_wire_out_253,
    output[1:0] io_V_wire_out_252,
    output[1:0] io_V_wire_out_251,
    output[1:0] io_V_wire_out_250,
    output[1:0] io_V_wire_out_249,
    output[1:0] io_V_wire_out_248,
    output[1:0] io_V_wire_out_247,
    output[1:0] io_V_wire_out_246,
    output[1:0] io_V_wire_out_245,
    output[1:0] io_V_wire_out_244,
    output[1:0] io_V_wire_out_243,
    output[1:0] io_V_wire_out_242,
    output[1:0] io_V_wire_out_241,
    output[1:0] io_V_wire_out_240,
    output[1:0] io_V_wire_out_239,
    output[1:0] io_V_wire_out_238,
    output[1:0] io_V_wire_out_237,
    output[1:0] io_V_wire_out_236,
    output[1:0] io_V_wire_out_235,
    output[1:0] io_V_wire_out_234,
    output[1:0] io_V_wire_out_233,
    output[1:0] io_V_wire_out_232,
    output[1:0] io_V_wire_out_231,
    output[1:0] io_V_wire_out_230,
    output[1:0] io_V_wire_out_229,
    output[1:0] io_V_wire_out_228,
    output[1:0] io_V_wire_out_227,
    output[1:0] io_V_wire_out_226,
    output[1:0] io_V_wire_out_225,
    output[1:0] io_V_wire_out_224,
    output[1:0] io_V_wire_out_223,
    output[1:0] io_V_wire_out_222,
    output[1:0] io_V_wire_out_221,
    output[1:0] io_V_wire_out_220,
    output[1:0] io_V_wire_out_219,
    output[1:0] io_V_wire_out_218,
    output[1:0] io_V_wire_out_217,
    output[1:0] io_V_wire_out_216,
    output[1:0] io_V_wire_out_215,
    output[1:0] io_V_wire_out_214,
    output[1:0] io_V_wire_out_213,
    output[1:0] io_V_wire_out_212,
    output[1:0] io_V_wire_out_211,
    output[1:0] io_V_wire_out_210,
    output[1:0] io_V_wire_out_209,
    output[1:0] io_V_wire_out_208,
    output[1:0] io_V_wire_out_207,
    output[1:0] io_V_wire_out_206,
    output[1:0] io_V_wire_out_205,
    output[1:0] io_V_wire_out_204,
    output[1:0] io_V_wire_out_203,
    output[1:0] io_V_wire_out_202,
    output[1:0] io_V_wire_out_201,
    output[1:0] io_V_wire_out_200,
    output[1:0] io_V_wire_out_199,
    output[1:0] io_V_wire_out_198,
    output[1:0] io_V_wire_out_197,
    output[1:0] io_V_wire_out_196,
    output[1:0] io_V_wire_out_195,
    output[1:0] io_V_wire_out_194,
    output[1:0] io_V_wire_out_193,
    output[1:0] io_V_wire_out_192,
    output[1:0] io_V_wire_out_191,
    output[1:0] io_V_wire_out_190,
    output[1:0] io_V_wire_out_189,
    output[1:0] io_V_wire_out_188,
    output[1:0] io_V_wire_out_187,
    output[1:0] io_V_wire_out_186,
    output[1:0] io_V_wire_out_185,
    output[1:0] io_V_wire_out_184,
    output[1:0] io_V_wire_out_183,
    output[1:0] io_V_wire_out_182,
    output[1:0] io_V_wire_out_181,
    output[1:0] io_V_wire_out_180,
    output[1:0] io_V_wire_out_179,
    output[1:0] io_V_wire_out_178,
    output[1:0] io_V_wire_out_177,
    output[1:0] io_V_wire_out_176,
    output[1:0] io_V_wire_out_175,
    output[1:0] io_V_wire_out_174,
    output[1:0] io_V_wire_out_173,
    output[1:0] io_V_wire_out_172,
    output[1:0] io_V_wire_out_171,
    output[1:0] io_V_wire_out_170,
    output[1:0] io_V_wire_out_169,
    output[1:0] io_V_wire_out_168,
    output[1:0] io_V_wire_out_167,
    output[1:0] io_V_wire_out_166,
    output[1:0] io_V_wire_out_165,
    output[1:0] io_V_wire_out_164,
    output[1:0] io_V_wire_out_163,
    output[1:0] io_V_wire_out_162,
    output[1:0] io_V_wire_out_161,
    output[1:0] io_V_wire_out_160,
    output[1:0] io_V_wire_out_159,
    output[1:0] io_V_wire_out_158,
    output[1:0] io_V_wire_out_157,
    output[1:0] io_V_wire_out_156,
    output[1:0] io_V_wire_out_155,
    output[1:0] io_V_wire_out_154,
    output[1:0] io_V_wire_out_153,
    output[1:0] io_V_wire_out_152,
    output[1:0] io_V_wire_out_151,
    output[1:0] io_V_wire_out_150,
    output[1:0] io_V_wire_out_149,
    output[1:0] io_V_wire_out_148,
    output[1:0] io_V_wire_out_147,
    output[1:0] io_V_wire_out_146,
    output[1:0] io_V_wire_out_145,
    output[1:0] io_V_wire_out_144,
    output[1:0] io_V_wire_out_143,
    output[1:0] io_V_wire_out_142,
    output[1:0] io_V_wire_out_141,
    output[1:0] io_V_wire_out_140,
    output[1:0] io_V_wire_out_139,
    output[1:0] io_V_wire_out_138,
    output[1:0] io_V_wire_out_137,
    output[1:0] io_V_wire_out_136,
    output[1:0] io_V_wire_out_135,
    output[1:0] io_V_wire_out_134,
    output[1:0] io_V_wire_out_133,
    output[1:0] io_V_wire_out_132,
    output[1:0] io_V_wire_out_131,
    output[1:0] io_V_wire_out_130,
    output[1:0] io_V_wire_out_129,
    output[1:0] io_V_wire_out_128,
    output[1:0] io_V_wire_out_127,
    output[1:0] io_V_wire_out_126,
    output[1:0] io_V_wire_out_125,
    output[1:0] io_V_wire_out_124,
    output[1:0] io_V_wire_out_123,
    output[1:0] io_V_wire_out_122,
    output[1:0] io_V_wire_out_121,
    output[1:0] io_V_wire_out_120,
    output[1:0] io_V_wire_out_119,
    output[1:0] io_V_wire_out_118,
    output[1:0] io_V_wire_out_117,
    output[1:0] io_V_wire_out_116,
    output[1:0] io_V_wire_out_115,
    output[1:0] io_V_wire_out_114,
    output[1:0] io_V_wire_out_113,
    output[1:0] io_V_wire_out_112,
    output[1:0] io_V_wire_out_111,
    output[1:0] io_V_wire_out_110,
    output[1:0] io_V_wire_out_109,
    output[1:0] io_V_wire_out_108,
    output[1:0] io_V_wire_out_107,
    output[1:0] io_V_wire_out_106,
    output[1:0] io_V_wire_out_105,
    output[1:0] io_V_wire_out_104,
    output[1:0] io_V_wire_out_103,
    output[1:0] io_V_wire_out_102,
    output[1:0] io_V_wire_out_101,
    output[1:0] io_V_wire_out_100,
    output[1:0] io_V_wire_out_99,
    output[1:0] io_V_wire_out_98,
    output[1:0] io_V_wire_out_97,
    output[1:0] io_V_wire_out_96,
    output[1:0] io_V_wire_out_95,
    output[1:0] io_V_wire_out_94,
    output[1:0] io_V_wire_out_93,
    output[1:0] io_V_wire_out_92,
    output[1:0] io_V_wire_out_91,
    output[1:0] io_V_wire_out_90,
    output[1:0] io_V_wire_out_89,
    output[1:0] io_V_wire_out_88,
    output[1:0] io_V_wire_out_87,
    output[1:0] io_V_wire_out_86,
    output[1:0] io_V_wire_out_85,
    output[1:0] io_V_wire_out_84,
    output[1:0] io_V_wire_out_83,
    output[1:0] io_V_wire_out_82,
    output[1:0] io_V_wire_out_81,
    output[1:0] io_V_wire_out_80,
    output[1:0] io_V_wire_out_79,
    output[1:0] io_V_wire_out_78,
    output[1:0] io_V_wire_out_77,
    output[1:0] io_V_wire_out_76,
    output[1:0] io_V_wire_out_75,
    output[1:0] io_V_wire_out_74,
    output[1:0] io_V_wire_out_73,
    output[1:0] io_V_wire_out_72,
    output[1:0] io_V_wire_out_71,
    output[1:0] io_V_wire_out_70,
    output[1:0] io_V_wire_out_69,
    output[1:0] io_V_wire_out_68,
    output[1:0] io_V_wire_out_67,
    output[1:0] io_V_wire_out_66,
    output[1:0] io_V_wire_out_65,
    output[1:0] io_V_wire_out_64,
    output[1:0] io_V_wire_out_63,
    output[1:0] io_V_wire_out_62,
    output[1:0] io_V_wire_out_61,
    output[1:0] io_V_wire_out_60,
    output[1:0] io_V_wire_out_59,
    output[1:0] io_V_wire_out_58,
    output[1:0] io_V_wire_out_57,
    output[1:0] io_V_wire_out_56,
    output[1:0] io_V_wire_out_55,
    output[1:0] io_V_wire_out_54,
    output[1:0] io_V_wire_out_53,
    output[1:0] io_V_wire_out_52,
    output[1:0] io_V_wire_out_51,
    output[1:0] io_V_wire_out_50,
    output[1:0] io_V_wire_out_49,
    output[1:0] io_V_wire_out_48,
    output[1:0] io_V_wire_out_47,
    output[1:0] io_V_wire_out_46,
    output[1:0] io_V_wire_out_45,
    output[1:0] io_V_wire_out_44,
    output[1:0] io_V_wire_out_43,
    output[1:0] io_V_wire_out_42,
    output[1:0] io_V_wire_out_41,
    output[1:0] io_V_wire_out_40,
    output[1:0] io_V_wire_out_39,
    output[1:0] io_V_wire_out_38,
    output[1:0] io_V_wire_out_37,
    output[1:0] io_V_wire_out_36,
    output[1:0] io_V_wire_out_35,
    output[1:0] io_V_wire_out_34,
    output[1:0] io_V_wire_out_33,
    output[1:0] io_V_wire_out_32,
    output[1:0] io_V_wire_out_31,
    output[1:0] io_V_wire_out_30,
    output[1:0] io_V_wire_out_29,
    output[1:0] io_V_wire_out_28,
    output[1:0] io_V_wire_out_27,
    output[1:0] io_V_wire_out_26,
    output[1:0] io_V_wire_out_25,
    output[1:0] io_V_wire_out_24,
    output[1:0] io_V_wire_out_23,
    output[1:0] io_V_wire_out_22,
    output[1:0] io_V_wire_out_21,
    output[1:0] io_V_wire_out_20,
    output[1:0] io_V_wire_out_19,
    output[1:0] io_V_wire_out_18,
    output[1:0] io_V_wire_out_17,
    output[1:0] io_V_wire_out_16,
    output[1:0] io_V_wire_out_15,
    output[1:0] io_V_wire_out_14,
    output[1:0] io_V_wire_out_13,
    output[1:0] io_V_wire_out_12,
    output[1:0] io_V_wire_out_11,
    output[1:0] io_V_wire_out_10,
    output[1:0] io_V_wire_out_9,
    output[1:0] io_V_wire_out_8,
    output[1:0] io_V_wire_out_7,
    output[1:0] io_V_wire_out_6,
    output[1:0] io_V_wire_out_5,
    output[1:0] io_V_wire_out_4,
    output[1:0] io_V_wire_out_3,
    output[1:0] io_V_wire_out_2,
    output[1:0] io_V_wire_out_1,
    output[1:0] io_V_wire_out_0,
    output[15:0] io_V_wire_en_22,
    output[15:0] io_V_wire_en_21,
    output[15:0] io_V_wire_en_20,
    output[15:0] io_V_wire_en_19,
    output[15:0] io_V_wire_en_18,
    output[15:0] io_V_wire_en_17,
    output[15:0] io_V_wire_en_16,
    output[15:0] io_V_wire_en_15,
    output[15:0] io_V_wire_en_14,
    output[15:0] io_V_wire_en_13,
    output[15:0] io_V_wire_en_12,
    output[15:0] io_V_wire_en_11,
    output[15:0] io_V_wire_en_10,
    output[15:0] io_V_wire_en_9,
    output[15:0] io_V_wire_en_8,
    output[15:0] io_V_wire_en_7,
    output[15:0] io_V_wire_en_6,
    output[15:0] io_V_wire_en_5,
    output[15:0] io_V_wire_en_4,
    output[15:0] io_V_wire_en_3,
    output[15:0] io_V_wire_en_2,
    output[15:0] io_V_wire_en_1,
    output[15:0] io_V_wire_en_0,
    input [1:0] io_G_wire_above_3,
    input [1:0] io_G_wire_above_2,
    input [1:0] io_G_wire_above_1,
    input [1:0] io_G_wire_above_0,
    input [1:0] io_H_wire_above_32,
    input [1:0] io_H_wire_above_31,
    input [1:0] io_H_wire_above_30,
    input [1:0] io_H_wire_above_29,
    input [1:0] io_H_wire_above_28,
    input [1:0] io_H_wire_above_27,
    input [1:0] io_H_wire_above_26,
    input [1:0] io_H_wire_above_25,
    input [1:0] io_H_wire_above_24,
    input [1:0] io_H_wire_above_23,
    input [1:0] io_H_wire_above_22,
    input [1:0] io_H_wire_above_21,
    input [1:0] io_H_wire_above_20,
    input [1:0] io_H_wire_above_19,
    input [1:0] io_H_wire_above_18,
    input [1:0] io_H_wire_above_17,
    input [1:0] io_H_wire_above_16,
    input [1:0] io_H_wire_above_15,
    input [1:0] io_H_wire_above_14,
    input [1:0] io_H_wire_above_13,
    input [1:0] io_H_wire_above_12,
    input [1:0] io_H_wire_above_11,
    input [1:0] io_H_wire_above_10,
    input [1:0] io_H_wire_above_9,
    input [1:0] io_H_wire_above_8,
    input [1:0] io_H_wire_above_7,
    input [1:0] io_H_wire_above_6,
    input [1:0] io_H_wire_above_5,
    input [1:0] io_H_wire_above_4,
    input [1:0] io_H_wire_above_3,
    input [1:0] io_H_wire_above_2,
    input [1:0] io_H_wire_above_1,
    input [1:0] io_H_wire_above_0,
    input [1:0] io_mem_bus_in_23,
    input [1:0] io_mem_bus_in_22,
    input [1:0] io_mem_bus_in_21,
    input [1:0] io_mem_bus_in_20,
    input [1:0] io_mem_bus_in_19,
    input [1:0] io_mem_bus_in_18,
    input [1:0] io_mem_bus_in_17,
    input [1:0] io_mem_bus_in_16,
    input [1:0] io_mem_bus_in_15,
    input [1:0] io_mem_bus_in_14,
    input [1:0] io_mem_bus_in_13,
    input [1:0] io_mem_bus_in_12,
    input [1:0] io_mem_bus_in_11,
    input [1:0] io_mem_bus_in_10,
    input [1:0] io_mem_bus_in_9,
    input [1:0] io_mem_bus_in_8,
    input [1:0] io_mem_bus_in_7,
    input [1:0] io_mem_bus_in_6,
    input [1:0] io_mem_bus_in_5,
    input [1:0] io_mem_bus_in_4,
    input [1:0] io_mem_bus_in_3,
    input [1:0] io_mem_bus_in_2,
    input [1:0] io_mem_bus_in_1,
    input [1:0] io_mem_bus_in_0,
    input [1:0] io_H_out_above_22,
    input [1:0] io_H_out_above_21,
    input [1:0] io_H_out_above_20,
    input [1:0] io_H_out_above_19,
    input [1:0] io_H_out_above_18,
    input [1:0] io_H_out_above_17,
    input [1:0] io_H_out_above_16,
    input [1:0] io_H_out_above_15,
    input [1:0] io_H_out_above_14,
    input [1:0] io_H_out_above_13,
    input [1:0] io_H_out_above_12,
    input [1:0] io_H_out_above_11,
    input [1:0] io_H_out_above_10,
    input [1:0] io_H_out_above_9,
    input [1:0] io_H_out_above_8,
    input [1:0] io_H_out_above_7,
    input [1:0] io_H_out_above_6,
    input [1:0] io_H_out_above_5,
    input [1:0] io_H_out_above_4,
    input [1:0] io_H_out_above_3,
    input [1:0] io_H_out_above_2,
    input [1:0] io_H_out_above_1,
    input [1:0] io_H_out_above_0,
    output[1:0] io_H_out_22,
    output[1:0] io_H_out_21,
    output[1:0] io_H_out_20,
    output[1:0] io_H_out_19,
    output[1:0] io_H_out_18,
    output[1:0] io_H_out_17,
    output[1:0] io_H_out_16,
    output[1:0] io_H_out_15,
    output[1:0] io_H_out_14,
    output[1:0] io_H_out_13,
    output[1:0] io_H_out_12,
    output[1:0] io_H_out_11,
    output[1:0] io_H_out_10,
    output[1:0] io_H_out_9,
    output[1:0] io_H_out_8,
    output[1:0] io_H_out_7,
    output[1:0] io_H_out_6,
    output[1:0] io_H_out_5,
    output[1:0] io_H_out_4,
    output[1:0] io_H_out_3,
    output[1:0] io_H_out_2,
    output[1:0] io_H_out_1,
    output[1:0] io_H_out_0,
    output[1:0] io_G_wire_below_3,
    output[1:0] io_G_wire_below_2,
    output[1:0] io_G_wire_below_1,
    output[1:0] io_G_wire_below_0,
    output[1:0] io_H_wire_below_32,
    output[1:0] io_H_wire_below_31,
    output[1:0] io_H_wire_below_30,
    output[1:0] io_H_wire_below_29,
    output[1:0] io_H_wire_below_28,
    output[1:0] io_H_wire_below_27,
    output[1:0] io_H_wire_below_26,
    output[1:0] io_H_wire_below_25,
    output[1:0] io_H_wire_below_24,
    output[1:0] io_H_wire_below_23,
    output[1:0] io_H_wire_below_22,
    output[1:0] io_H_wire_below_21,
    output[1:0] io_H_wire_below_20,
    output[1:0] io_H_wire_below_19,
    output[1:0] io_H_wire_below_18,
    output[1:0] io_H_wire_below_17,
    output[1:0] io_H_wire_below_16,
    output[1:0] io_H_wire_below_15,
    output[1:0] io_H_wire_below_14,
    output[1:0] io_H_wire_below_13,
    output[1:0] io_H_wire_below_12,
    output[1:0] io_H_wire_below_11,
    output[1:0] io_H_wire_below_10,
    output[1:0] io_H_wire_below_9,
    output[1:0] io_H_wire_below_8,
    output[1:0] io_H_wire_below_7,
    output[1:0] io_H_wire_below_6,
    output[1:0] io_H_wire_below_5,
    output[1:0] io_H_wire_below_4,
    output[1:0] io_H_wire_below_3,
    output[1:0] io_H_wire_below_2,
    output[1:0] io_H_wire_below_1,
    output[1:0] io_H_wire_below_0,
    input  io_row_en,
    input  io_config_or_load,
    input  io_D_or_Z,
    output[1:0] io_mem_bus_out_23,
    output[1:0] io_mem_bus_out_22,
    output[1:0] io_mem_bus_out_21,
    output[1:0] io_mem_bus_out_20,
    output[1:0] io_mem_bus_out_19,
    output[1:0] io_mem_bus_out_18,
    output[1:0] io_mem_bus_out_17,
    output[1:0] io_mem_bus_out_16,
    output[1:0] io_mem_bus_out_15,
    output[1:0] io_mem_bus_out_14,
    output[1:0] io_mem_bus_out_13,
    output[1:0] io_mem_bus_out_12,
    output[1:0] io_mem_bus_out_11,
    output[1:0] io_mem_bus_out_10,
    output[1:0] io_mem_bus_out_9,
    output[1:0] io_mem_bus_out_8,
    output[1:0] io_mem_bus_out_7,
    output[1:0] io_mem_bus_out_6,
    output[1:0] io_mem_bus_out_5,
    output[1:0] io_mem_bus_out_4,
    output[1:0] io_mem_bus_out_3,
    output[1:0] io_mem_bus_out_2,
    output[1:0] io_mem_bus_out_1,
    output[1:0] io_mem_bus_out_0
);

  wire[1:0] T0;
  wire T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire[1:0] T28;
  wire[1:0] T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire[1:0] T42;
  wire[1:0] T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire[1:0] T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire[1:0] T50;
  wire[1:0] T51;
  wire[1:0] T52;
  wire[1:0] T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire[1:0] T60;
  wire[1:0] T61;
  wire[1:0] T62;
  wire[1:0] T63;
  wire[1:0] T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire[1:0] T70;
  wire[1:0] T71;
  wire[22:0] G_wire_below_en_3;
  wire[22:0] T5018;
  wire[23:0] T72;
  wire[23:0] T5019;
  wire[22:0] T73;
  wire[22:0] T5020;
  wire[21:0] T74;
  wire[21:0] T5021;
  wire[20:0] T75;
  wire[20:0] T5022;
  wire[19:0] T76;
  wire[19:0] T5023;
  wire[18:0] T77;
  wire[18:0] T5024;
  wire[17:0] T78;
  wire[17:0] T5025;
  wire[16:0] T79;
  wire[16:0] T5026;
  wire[15:0] T80;
  wire[15:0] T5027;
  wire[14:0] T81;
  wire[14:0] T5028;
  wire[13:0] T82;
  wire[13:0] T5029;
  wire[12:0] T83;
  wire[12:0] T5030;
  wire[11:0] T84;
  wire[11:0] T5031;
  wire[10:0] T85;
  wire[10:0] T5032;
  wire[9:0] T86;
  wire[9:0] T5033;
  wire[8:0] T87;
  wire[8:0] T5034;
  wire[7:0] T88;
  wire[7:0] T5035;
  wire[6:0] T89;
  wire[6:0] T5036;
  wire[5:0] T90;
  wire[5:0] T5037;
  wire[4:0] T91;
  wire[4:0] T5038;
  wire[3:0] T92;
  wire[3:0] T5039;
  wire[2:0] T93;
  wire[2:0] T5040;
  wire[1:0] T94;
  wire[1:0] T95;
  wire[1:0] T96;
  wire[1:0] T97;
  wire[1:0] T5041;
  wire T98;
  wire T99;
  wire[1:0] T100;
  wire[1:0] T101;
  wire T102;
  wire T103;
  wire[1:0] T104;
  wire T105;
  wire T106;
  wire[2:0] T107;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] T5042;
  wire T110;
  wire T111;
  wire[2:0] T112;
  wire[2:0] T113;
  wire[2:0] T5043;
  wire T114;
  wire T115;
  wire[1:0] T116;
  wire T117;
  wire T118;
  wire[3:0] T119;
  wire[3:0] T120;
  wire[3:0] T121;
  wire[3:0] T5044;
  wire T122;
  wire T123;
  wire[3:0] T124;
  wire[3:0] T125;
  wire[3:0] T5045;
  wire T126;
  wire T127;
  wire[1:0] T128;
  wire T129;
  wire T130;
  wire[4:0] T131;
  wire[4:0] T132;
  wire[4:0] T133;
  wire[4:0] T5046;
  wire T134;
  wire T135;
  wire[4:0] T136;
  wire[4:0] T137;
  wire[4:0] T5047;
  wire T138;
  wire T139;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire[5:0] T143;
  wire[5:0] T144;
  wire[5:0] T145;
  wire[5:0] T5048;
  wire T146;
  wire T147;
  wire[5:0] T148;
  wire[5:0] T149;
  wire[5:0] T5049;
  wire T150;
  wire T151;
  wire[1:0] T152;
  wire T153;
  wire T154;
  wire[6:0] T155;
  wire[6:0] T156;
  wire[6:0] T157;
  wire[6:0] T5050;
  wire T158;
  wire T159;
  wire[6:0] T160;
  wire[6:0] T161;
  wire[6:0] T5051;
  wire T162;
  wire T163;
  wire[1:0] T164;
  wire T165;
  wire T166;
  wire[7:0] T167;
  wire[7:0] T168;
  wire[7:0] T169;
  wire[7:0] T5052;
  wire T170;
  wire T171;
  wire[7:0] T172;
  wire[7:0] T173;
  wire[7:0] T5053;
  wire T174;
  wire T175;
  wire[1:0] T176;
  wire T177;
  wire T178;
  wire[8:0] T179;
  wire[8:0] T180;
  wire[8:0] T181;
  wire[8:0] T5054;
  wire T182;
  wire T183;
  wire[8:0] T184;
  wire[8:0] T185;
  wire[8:0] T5055;
  wire T186;
  wire T187;
  wire[1:0] T188;
  wire T189;
  wire T190;
  wire[9:0] T191;
  wire[9:0] T192;
  wire[9:0] T193;
  wire[9:0] T5056;
  wire T194;
  wire T195;
  wire[9:0] T196;
  wire[9:0] T197;
  wire[9:0] T5057;
  wire T198;
  wire T199;
  wire[1:0] T200;
  wire T201;
  wire T202;
  wire[10:0] T203;
  wire[10:0] T204;
  wire[10:0] T205;
  wire[10:0] T5058;
  wire T206;
  wire T207;
  wire[10:0] T208;
  wire[10:0] T209;
  wire[10:0] T5059;
  wire T210;
  wire T211;
  wire[1:0] T212;
  wire T213;
  wire T214;
  wire[11:0] T215;
  wire[11:0] T216;
  wire[11:0] T217;
  wire[11:0] T5060;
  wire T218;
  wire T219;
  wire[11:0] T220;
  wire[11:0] T221;
  wire[11:0] T5061;
  wire T222;
  wire T223;
  wire[1:0] T224;
  wire T225;
  wire T226;
  wire[12:0] T227;
  wire[12:0] T228;
  wire[12:0] T229;
  wire[12:0] T5062;
  wire T230;
  wire T231;
  wire[12:0] T232;
  wire[12:0] T233;
  wire[12:0] T5063;
  wire T234;
  wire T235;
  wire[1:0] T236;
  wire T237;
  wire T238;
  wire[13:0] T239;
  wire[13:0] T240;
  wire[13:0] T241;
  wire[13:0] T5064;
  wire T242;
  wire T243;
  wire[13:0] T244;
  wire[13:0] T245;
  wire[13:0] T5065;
  wire T246;
  wire T247;
  wire[1:0] T248;
  wire T249;
  wire T250;
  wire[14:0] T251;
  wire[14:0] T252;
  wire[14:0] T253;
  wire[14:0] T5066;
  wire T254;
  wire T255;
  wire[14:0] T256;
  wire[14:0] T257;
  wire[14:0] T5067;
  wire T258;
  wire T259;
  wire[1:0] T260;
  wire T261;
  wire T262;
  wire[15:0] T263;
  wire[15:0] T264;
  wire[15:0] T265;
  wire[15:0] T5068;
  wire T266;
  wire T267;
  wire[15:0] T268;
  wire[15:0] T269;
  wire[15:0] T5069;
  wire T270;
  wire T271;
  wire[1:0] T272;
  wire T273;
  wire T274;
  wire[16:0] T275;
  wire[16:0] T276;
  wire[16:0] T277;
  wire[16:0] T5070;
  wire T278;
  wire T279;
  wire[16:0] T280;
  wire[16:0] T281;
  wire[16:0] T5071;
  wire T282;
  wire T283;
  wire[1:0] T284;
  wire T285;
  wire T286;
  wire[17:0] T287;
  wire[17:0] T288;
  wire[17:0] T289;
  wire[17:0] T5072;
  wire T290;
  wire T291;
  wire[17:0] T292;
  wire[17:0] T293;
  wire[17:0] T5073;
  wire T294;
  wire T295;
  wire[1:0] T296;
  wire T297;
  wire T298;
  wire[18:0] T299;
  wire[18:0] T300;
  wire[18:0] T301;
  wire[18:0] T5074;
  wire T302;
  wire T303;
  wire[18:0] T304;
  wire[18:0] T305;
  wire[18:0] T5075;
  wire T306;
  wire T307;
  wire[1:0] T308;
  wire T309;
  wire T310;
  wire[19:0] T311;
  wire[19:0] T312;
  wire[19:0] T313;
  wire[19:0] T5076;
  wire T314;
  wire T315;
  wire[19:0] T316;
  wire[19:0] T317;
  wire[19:0] T5077;
  wire T318;
  wire T319;
  wire[1:0] T320;
  wire T321;
  wire T322;
  wire[20:0] T323;
  wire[20:0] T324;
  wire[20:0] T325;
  wire[20:0] T5078;
  wire T326;
  wire T327;
  wire[20:0] T328;
  wire[20:0] T329;
  wire[20:0] T5079;
  wire T330;
  wire T331;
  wire[1:0] T332;
  wire T333;
  wire T334;
  wire[21:0] T335;
  wire[21:0] T336;
  wire[21:0] T337;
  wire[21:0] T5080;
  wire T338;
  wire T339;
  wire[21:0] T340;
  wire[21:0] T341;
  wire[21:0] T5081;
  wire T342;
  wire T343;
  wire[1:0] T344;
  wire T345;
  wire T346;
  wire[22:0] T347;
  wire[22:0] T348;
  wire[22:0] T349;
  wire[22:0] T5082;
  wire T350;
  wire T351;
  wire[22:0] T352;
  wire[22:0] T353;
  wire[22:0] T5083;
  wire T354;
  wire T355;
  wire[1:0] T356;
  wire T357;
  wire T358;
  wire[23:0] T359;
  wire[23:0] T360;
  wire[23:0] T361;
  wire[23:0] T5084;
  wire T362;
  wire T363;
  wire[23:0] T364;
  wire[23:0] T365;
  wire[23:0] T5085;
  wire T366;
  wire T367;
  wire[1:0] T368;
  wire T369;
  wire T370;
  wire[1:0] G_wire_outs_0;
  wire[1:0] G_wire_outs_1;
  wire[1:0] G_wire_outs_2;
  wire[1:0] G_wire_outs_3;
  wire[1:0] G_wire_outs_4;
  wire[1:0] G_wire_outs_5;
  wire[1:0] G_wire_outs_6;
  wire[1:0] G_wire_outs_7;
  wire[1:0] G_wire_outs_8;
  wire[1:0] G_wire_outs_9;
  wire[1:0] G_wire_outs_10;
  wire[1:0] G_wire_outs_11;
  wire[1:0] G_wire_outs_12;
  wire[1:0] G_wire_outs_13;
  wire[1:0] G_wire_outs_14;
  wire[1:0] G_wire_outs_15;
  wire[1:0] G_wire_outs_16;
  wire[1:0] G_wire_outs_17;
  wire[1:0] G_wire_outs_18;
  wire[1:0] G_wire_outs_19;
  wire[1:0] G_wire_outs_20;
  wire[1:0] G_wire_outs_21;
  wire[1:0] G_wire_outs_22;
  wire[22:0] G_wire_below_en_2;
  wire[22:0] T5086;
  wire[23:0] T371;
  wire[23:0] T5087;
  wire[22:0] T372;
  wire[22:0] T5088;
  wire[21:0] T373;
  wire[21:0] T5089;
  wire[20:0] T374;
  wire[20:0] T5090;
  wire[19:0] T375;
  wire[19:0] T5091;
  wire[18:0] T376;
  wire[18:0] T5092;
  wire[17:0] T377;
  wire[17:0] T5093;
  wire[16:0] T378;
  wire[16:0] T5094;
  wire[15:0] T379;
  wire[15:0] T5095;
  wire[14:0] T380;
  wire[14:0] T5096;
  wire[13:0] T381;
  wire[13:0] T5097;
  wire[12:0] T382;
  wire[12:0] T5098;
  wire[11:0] T383;
  wire[11:0] T5099;
  wire[10:0] T384;
  wire[10:0] T5100;
  wire[9:0] T385;
  wire[9:0] T5101;
  wire[8:0] T386;
  wire[8:0] T5102;
  wire[7:0] T387;
  wire[7:0] T5103;
  wire[6:0] T388;
  wire[6:0] T5104;
  wire[5:0] T389;
  wire[5:0] T5105;
  wire[4:0] T390;
  wire[4:0] T5106;
  wire[3:0] T391;
  wire[3:0] T5107;
  wire[2:0] T392;
  wire[2:0] T5108;
  wire[1:0] T393;
  wire[1:0] T394;
  wire[1:0] T395;
  wire[1:0] T396;
  wire[1:0] T5109;
  wire T397;
  wire T398;
  wire[1:0] T399;
  wire[1:0] T400;
  wire T401;
  wire T402;
  wire[2:0] T403;
  wire[2:0] T404;
  wire[2:0] T405;
  wire[2:0] T5110;
  wire T406;
  wire T407;
  wire[2:0] T408;
  wire[2:0] T409;
  wire[2:0] T5111;
  wire T410;
  wire T411;
  wire[3:0] T412;
  wire[3:0] T413;
  wire[3:0] T414;
  wire[3:0] T5112;
  wire T415;
  wire T416;
  wire[3:0] T417;
  wire[3:0] T418;
  wire[3:0] T5113;
  wire T419;
  wire T420;
  wire[4:0] T421;
  wire[4:0] T422;
  wire[4:0] T423;
  wire[4:0] T5114;
  wire T424;
  wire T425;
  wire[4:0] T426;
  wire[4:0] T427;
  wire[4:0] T5115;
  wire T428;
  wire T429;
  wire[5:0] T430;
  wire[5:0] T431;
  wire[5:0] T432;
  wire[5:0] T5116;
  wire T433;
  wire T434;
  wire[5:0] T435;
  wire[5:0] T436;
  wire[5:0] T5117;
  wire T437;
  wire T438;
  wire[6:0] T439;
  wire[6:0] T440;
  wire[6:0] T441;
  wire[6:0] T5118;
  wire T442;
  wire T443;
  wire[6:0] T444;
  wire[6:0] T445;
  wire[6:0] T5119;
  wire T446;
  wire T447;
  wire[7:0] T448;
  wire[7:0] T449;
  wire[7:0] T450;
  wire[7:0] T5120;
  wire T451;
  wire T452;
  wire[7:0] T453;
  wire[7:0] T454;
  wire[7:0] T5121;
  wire T455;
  wire T456;
  wire[8:0] T457;
  wire[8:0] T458;
  wire[8:0] T459;
  wire[8:0] T5122;
  wire T460;
  wire T461;
  wire[8:0] T462;
  wire[8:0] T463;
  wire[8:0] T5123;
  wire T464;
  wire T465;
  wire[9:0] T466;
  wire[9:0] T467;
  wire[9:0] T468;
  wire[9:0] T5124;
  wire T469;
  wire T470;
  wire[9:0] T471;
  wire[9:0] T472;
  wire[9:0] T5125;
  wire T473;
  wire T474;
  wire[10:0] T475;
  wire[10:0] T476;
  wire[10:0] T477;
  wire[10:0] T5126;
  wire T478;
  wire T479;
  wire[10:0] T480;
  wire[10:0] T481;
  wire[10:0] T5127;
  wire T482;
  wire T483;
  wire[11:0] T484;
  wire[11:0] T485;
  wire[11:0] T486;
  wire[11:0] T5128;
  wire T487;
  wire T488;
  wire[11:0] T489;
  wire[11:0] T490;
  wire[11:0] T5129;
  wire T491;
  wire T492;
  wire[12:0] T493;
  wire[12:0] T494;
  wire[12:0] T495;
  wire[12:0] T5130;
  wire T496;
  wire T497;
  wire[12:0] T498;
  wire[12:0] T499;
  wire[12:0] T5131;
  wire T500;
  wire T501;
  wire[13:0] T502;
  wire[13:0] T503;
  wire[13:0] T504;
  wire[13:0] T5132;
  wire T505;
  wire T506;
  wire[13:0] T507;
  wire[13:0] T508;
  wire[13:0] T5133;
  wire T509;
  wire T510;
  wire[14:0] T511;
  wire[14:0] T512;
  wire[14:0] T513;
  wire[14:0] T5134;
  wire T514;
  wire T515;
  wire[14:0] T516;
  wire[14:0] T517;
  wire[14:0] T5135;
  wire T518;
  wire T519;
  wire[15:0] T520;
  wire[15:0] T521;
  wire[15:0] T522;
  wire[15:0] T5136;
  wire T523;
  wire T524;
  wire[15:0] T525;
  wire[15:0] T526;
  wire[15:0] T5137;
  wire T527;
  wire T528;
  wire[16:0] T529;
  wire[16:0] T530;
  wire[16:0] T531;
  wire[16:0] T5138;
  wire T532;
  wire T533;
  wire[16:0] T534;
  wire[16:0] T535;
  wire[16:0] T5139;
  wire T536;
  wire T537;
  wire[17:0] T538;
  wire[17:0] T539;
  wire[17:0] T540;
  wire[17:0] T5140;
  wire T541;
  wire T542;
  wire[17:0] T543;
  wire[17:0] T544;
  wire[17:0] T5141;
  wire T545;
  wire T546;
  wire[18:0] T547;
  wire[18:0] T548;
  wire[18:0] T549;
  wire[18:0] T5142;
  wire T550;
  wire T551;
  wire[18:0] T552;
  wire[18:0] T553;
  wire[18:0] T5143;
  wire T554;
  wire T555;
  wire[19:0] T556;
  wire[19:0] T557;
  wire[19:0] T558;
  wire[19:0] T5144;
  wire T559;
  wire T560;
  wire[19:0] T561;
  wire[19:0] T562;
  wire[19:0] T5145;
  wire T563;
  wire T564;
  wire[20:0] T565;
  wire[20:0] T566;
  wire[20:0] T567;
  wire[20:0] T5146;
  wire T568;
  wire T569;
  wire[20:0] T570;
  wire[20:0] T571;
  wire[20:0] T5147;
  wire T572;
  wire T573;
  wire[21:0] T574;
  wire[21:0] T575;
  wire[21:0] T576;
  wire[21:0] T5148;
  wire T577;
  wire T578;
  wire[21:0] T579;
  wire[21:0] T580;
  wire[21:0] T5149;
  wire T581;
  wire T582;
  wire[22:0] T583;
  wire[22:0] T584;
  wire[22:0] T585;
  wire[22:0] T5150;
  wire T586;
  wire T587;
  wire[22:0] T588;
  wire[22:0] T589;
  wire[22:0] T5151;
  wire T590;
  wire T591;
  wire[23:0] T592;
  wire[23:0] T593;
  wire[23:0] T594;
  wire[23:0] T5152;
  wire T595;
  wire T596;
  wire[23:0] T597;
  wire[23:0] T598;
  wire[23:0] T5153;
  wire T599;
  wire T600;
  wire[22:0] G_wire_below_en_1;
  wire[22:0] T5154;
  wire[23:0] T601;
  wire[23:0] T5155;
  wire[22:0] T602;
  wire[22:0] T5156;
  wire[21:0] T603;
  wire[21:0] T5157;
  wire[20:0] T604;
  wire[20:0] T5158;
  wire[19:0] T605;
  wire[19:0] T5159;
  wire[18:0] T606;
  wire[18:0] T5160;
  wire[17:0] T607;
  wire[17:0] T5161;
  wire[16:0] T608;
  wire[16:0] T5162;
  wire[15:0] T609;
  wire[15:0] T5163;
  wire[14:0] T610;
  wire[14:0] T5164;
  wire[13:0] T611;
  wire[13:0] T5165;
  wire[12:0] T612;
  wire[12:0] T5166;
  wire[11:0] T613;
  wire[11:0] T5167;
  wire[10:0] T614;
  wire[10:0] T5168;
  wire[9:0] T615;
  wire[9:0] T5169;
  wire[8:0] T616;
  wire[8:0] T5170;
  wire[7:0] T617;
  wire[7:0] T5171;
  wire[6:0] T618;
  wire[6:0] T5172;
  wire[5:0] T619;
  wire[5:0] T5173;
  wire[4:0] T620;
  wire[4:0] T5174;
  wire[3:0] T621;
  wire[3:0] T5175;
  wire[2:0] T622;
  wire[2:0] T5176;
  wire[1:0] T623;
  wire[1:0] T624;
  wire[1:0] T625;
  wire[1:0] T626;
  wire[1:0] T5177;
  wire T627;
  wire T628;
  wire[1:0] T629;
  wire[1:0] T630;
  wire T631;
  wire T632;
  wire[2:0] T633;
  wire[2:0] T634;
  wire[2:0] T635;
  wire[2:0] T5178;
  wire T636;
  wire T637;
  wire[2:0] T638;
  wire[2:0] T639;
  wire[2:0] T5179;
  wire T640;
  wire T641;
  wire[3:0] T642;
  wire[3:0] T643;
  wire[3:0] T644;
  wire[3:0] T5180;
  wire T645;
  wire T646;
  wire[3:0] T647;
  wire[3:0] T648;
  wire[3:0] T5181;
  wire T649;
  wire T650;
  wire[4:0] T651;
  wire[4:0] T652;
  wire[4:0] T653;
  wire[4:0] T5182;
  wire T654;
  wire T655;
  wire[4:0] T656;
  wire[4:0] T657;
  wire[4:0] T5183;
  wire T658;
  wire T659;
  wire[5:0] T660;
  wire[5:0] T661;
  wire[5:0] T662;
  wire[5:0] T5184;
  wire T663;
  wire T664;
  wire[5:0] T665;
  wire[5:0] T666;
  wire[5:0] T5185;
  wire T667;
  wire T668;
  wire[6:0] T669;
  wire[6:0] T670;
  wire[6:0] T671;
  wire[6:0] T5186;
  wire T672;
  wire T673;
  wire[6:0] T674;
  wire[6:0] T675;
  wire[6:0] T5187;
  wire T676;
  wire T677;
  wire[7:0] T678;
  wire[7:0] T679;
  wire[7:0] T680;
  wire[7:0] T5188;
  wire T681;
  wire T682;
  wire[7:0] T683;
  wire[7:0] T684;
  wire[7:0] T5189;
  wire T685;
  wire T686;
  wire[8:0] T687;
  wire[8:0] T688;
  wire[8:0] T689;
  wire[8:0] T5190;
  wire T690;
  wire T691;
  wire[8:0] T692;
  wire[8:0] T693;
  wire[8:0] T5191;
  wire T694;
  wire T695;
  wire[9:0] T696;
  wire[9:0] T697;
  wire[9:0] T698;
  wire[9:0] T5192;
  wire T699;
  wire T700;
  wire[9:0] T701;
  wire[9:0] T702;
  wire[9:0] T5193;
  wire T703;
  wire T704;
  wire[10:0] T705;
  wire[10:0] T706;
  wire[10:0] T707;
  wire[10:0] T5194;
  wire T708;
  wire T709;
  wire[10:0] T710;
  wire[10:0] T711;
  wire[10:0] T5195;
  wire T712;
  wire T713;
  wire[11:0] T714;
  wire[11:0] T715;
  wire[11:0] T716;
  wire[11:0] T5196;
  wire T717;
  wire T718;
  wire[11:0] T719;
  wire[11:0] T720;
  wire[11:0] T5197;
  wire T721;
  wire T722;
  wire[12:0] T723;
  wire[12:0] T724;
  wire[12:0] T725;
  wire[12:0] T5198;
  wire T726;
  wire T727;
  wire[12:0] T728;
  wire[12:0] T729;
  wire[12:0] T5199;
  wire T730;
  wire T731;
  wire[13:0] T732;
  wire[13:0] T733;
  wire[13:0] T734;
  wire[13:0] T5200;
  wire T735;
  wire T736;
  wire[13:0] T737;
  wire[13:0] T738;
  wire[13:0] T5201;
  wire T739;
  wire T740;
  wire[14:0] T741;
  wire[14:0] T742;
  wire[14:0] T743;
  wire[14:0] T5202;
  wire T744;
  wire T745;
  wire[14:0] T746;
  wire[14:0] T747;
  wire[14:0] T5203;
  wire T748;
  wire T749;
  wire[15:0] T750;
  wire[15:0] T751;
  wire[15:0] T752;
  wire[15:0] T5204;
  wire T753;
  wire T754;
  wire[15:0] T755;
  wire[15:0] T756;
  wire[15:0] T5205;
  wire T757;
  wire T758;
  wire[16:0] T759;
  wire[16:0] T760;
  wire[16:0] T761;
  wire[16:0] T5206;
  wire T762;
  wire T763;
  wire[16:0] T764;
  wire[16:0] T765;
  wire[16:0] T5207;
  wire T766;
  wire T767;
  wire[17:0] T768;
  wire[17:0] T769;
  wire[17:0] T770;
  wire[17:0] T5208;
  wire T771;
  wire T772;
  wire[17:0] T773;
  wire[17:0] T774;
  wire[17:0] T5209;
  wire T775;
  wire T776;
  wire[18:0] T777;
  wire[18:0] T778;
  wire[18:0] T779;
  wire[18:0] T5210;
  wire T780;
  wire T781;
  wire[18:0] T782;
  wire[18:0] T783;
  wire[18:0] T5211;
  wire T784;
  wire T785;
  wire[19:0] T786;
  wire[19:0] T787;
  wire[19:0] T788;
  wire[19:0] T5212;
  wire T789;
  wire T790;
  wire[19:0] T791;
  wire[19:0] T792;
  wire[19:0] T5213;
  wire T793;
  wire T794;
  wire[20:0] T795;
  wire[20:0] T796;
  wire[20:0] T797;
  wire[20:0] T5214;
  wire T798;
  wire T799;
  wire[20:0] T800;
  wire[20:0] T801;
  wire[20:0] T5215;
  wire T802;
  wire T803;
  wire[21:0] T804;
  wire[21:0] T805;
  wire[21:0] T806;
  wire[21:0] T5216;
  wire T807;
  wire T808;
  wire[21:0] T809;
  wire[21:0] T810;
  wire[21:0] T5217;
  wire T811;
  wire T812;
  wire[22:0] T813;
  wire[22:0] T814;
  wire[22:0] T815;
  wire[22:0] T5218;
  wire T816;
  wire T817;
  wire[22:0] T818;
  wire[22:0] T819;
  wire[22:0] T5219;
  wire T820;
  wire T821;
  wire[23:0] T822;
  wire[23:0] T823;
  wire[23:0] T824;
  wire[23:0] T5220;
  wire T825;
  wire T826;
  wire[23:0] T827;
  wire[23:0] T828;
  wire[23:0] T5221;
  wire T829;
  wire T830;
  wire[22:0] G_wire_below_en_0;
  wire[22:0] T5222;
  wire[23:0] T831;
  wire[23:0] T5223;
  wire[22:0] T832;
  wire[22:0] T5224;
  wire[21:0] T833;
  wire[21:0] T5225;
  wire[20:0] T834;
  wire[20:0] T5226;
  wire[19:0] T835;
  wire[19:0] T5227;
  wire[18:0] T836;
  wire[18:0] T5228;
  wire[17:0] T837;
  wire[17:0] T5229;
  wire[16:0] T838;
  wire[16:0] T5230;
  wire[15:0] T839;
  wire[15:0] T5231;
  wire[14:0] T840;
  wire[14:0] T5232;
  wire[13:0] T841;
  wire[13:0] T5233;
  wire[12:0] T842;
  wire[12:0] T5234;
  wire[11:0] T843;
  wire[11:0] T5235;
  wire[10:0] T844;
  wire[10:0] T5236;
  wire[9:0] T845;
  wire[9:0] T5237;
  wire[8:0] T846;
  wire[8:0] T5238;
  wire[7:0] T847;
  wire[7:0] T5239;
  wire[6:0] T848;
  wire[6:0] T5240;
  wire[5:0] T849;
  wire[5:0] T5241;
  wire[4:0] T850;
  wire[4:0] T5242;
  wire[3:0] T851;
  wire[3:0] T5243;
  wire[2:0] T852;
  wire[2:0] T5244;
  wire[1:0] T853;
  wire[1:0] T854;
  wire[1:0] T855;
  wire[1:0] T856;
  wire[1:0] T5245;
  wire T857;
  wire T858;
  wire[1:0] T859;
  wire[1:0] T860;
  wire T861;
  wire T862;
  wire[2:0] T863;
  wire[2:0] T864;
  wire[2:0] T865;
  wire[2:0] T5246;
  wire T866;
  wire T867;
  wire[2:0] T868;
  wire[2:0] T869;
  wire[2:0] T5247;
  wire T870;
  wire T871;
  wire[3:0] T872;
  wire[3:0] T873;
  wire[3:0] T874;
  wire[3:0] T5248;
  wire T875;
  wire T876;
  wire[3:0] T877;
  wire[3:0] T878;
  wire[3:0] T5249;
  wire T879;
  wire T880;
  wire[4:0] T881;
  wire[4:0] T882;
  wire[4:0] T883;
  wire[4:0] T5250;
  wire T884;
  wire T885;
  wire[4:0] T886;
  wire[4:0] T887;
  wire[4:0] T5251;
  wire T888;
  wire T889;
  wire[5:0] T890;
  wire[5:0] T891;
  wire[5:0] T892;
  wire[5:0] T5252;
  wire T893;
  wire T894;
  wire[5:0] T895;
  wire[5:0] T896;
  wire[5:0] T5253;
  wire T897;
  wire T898;
  wire[6:0] T899;
  wire[6:0] T900;
  wire[6:0] T901;
  wire[6:0] T5254;
  wire T902;
  wire T903;
  wire[6:0] T904;
  wire[6:0] T905;
  wire[6:0] T5255;
  wire T906;
  wire T907;
  wire[7:0] T908;
  wire[7:0] T909;
  wire[7:0] T910;
  wire[7:0] T5256;
  wire T911;
  wire T912;
  wire[7:0] T913;
  wire[7:0] T914;
  wire[7:0] T5257;
  wire T915;
  wire T916;
  wire[8:0] T917;
  wire[8:0] T918;
  wire[8:0] T919;
  wire[8:0] T5258;
  wire T920;
  wire T921;
  wire[8:0] T922;
  wire[8:0] T923;
  wire[8:0] T5259;
  wire T924;
  wire T925;
  wire[9:0] T926;
  wire[9:0] T927;
  wire[9:0] T928;
  wire[9:0] T5260;
  wire T929;
  wire T930;
  wire[9:0] T931;
  wire[9:0] T932;
  wire[9:0] T5261;
  wire T933;
  wire T934;
  wire[10:0] T935;
  wire[10:0] T936;
  wire[10:0] T937;
  wire[10:0] T5262;
  wire T938;
  wire T939;
  wire[10:0] T940;
  wire[10:0] T941;
  wire[10:0] T5263;
  wire T942;
  wire T943;
  wire[11:0] T944;
  wire[11:0] T945;
  wire[11:0] T946;
  wire[11:0] T5264;
  wire T947;
  wire T948;
  wire[11:0] T949;
  wire[11:0] T950;
  wire[11:0] T5265;
  wire T951;
  wire T952;
  wire[12:0] T953;
  wire[12:0] T954;
  wire[12:0] T955;
  wire[12:0] T5266;
  wire T956;
  wire T957;
  wire[12:0] T958;
  wire[12:0] T959;
  wire[12:0] T5267;
  wire T960;
  wire T961;
  wire[13:0] T962;
  wire[13:0] T963;
  wire[13:0] T964;
  wire[13:0] T5268;
  wire T965;
  wire T966;
  wire[13:0] T967;
  wire[13:0] T968;
  wire[13:0] T5269;
  wire T969;
  wire T970;
  wire[14:0] T971;
  wire[14:0] T972;
  wire[14:0] T973;
  wire[14:0] T5270;
  wire T974;
  wire T975;
  wire[14:0] T976;
  wire[14:0] T977;
  wire[14:0] T5271;
  wire T978;
  wire T979;
  wire[15:0] T980;
  wire[15:0] T981;
  wire[15:0] T982;
  wire[15:0] T5272;
  wire T983;
  wire T984;
  wire[15:0] T985;
  wire[15:0] T986;
  wire[15:0] T5273;
  wire T987;
  wire T988;
  wire[16:0] T989;
  wire[16:0] T990;
  wire[16:0] T991;
  wire[16:0] T5274;
  wire T992;
  wire T993;
  wire[16:0] T994;
  wire[16:0] T995;
  wire[16:0] T5275;
  wire T996;
  wire T997;
  wire[17:0] T998;
  wire[17:0] T999;
  wire[17:0] T1000;
  wire[17:0] T5276;
  wire T1001;
  wire T1002;
  wire[17:0] T1003;
  wire[17:0] T1004;
  wire[17:0] T5277;
  wire T1005;
  wire T1006;
  wire[18:0] T1007;
  wire[18:0] T1008;
  wire[18:0] T1009;
  wire[18:0] T5278;
  wire T1010;
  wire T1011;
  wire[18:0] T1012;
  wire[18:0] T1013;
  wire[18:0] T5279;
  wire T1014;
  wire T1015;
  wire[19:0] T1016;
  wire[19:0] T1017;
  wire[19:0] T1018;
  wire[19:0] T5280;
  wire T1019;
  wire T1020;
  wire[19:0] T1021;
  wire[19:0] T1022;
  wire[19:0] T5281;
  wire T1023;
  wire T1024;
  wire[20:0] T1025;
  wire[20:0] T1026;
  wire[20:0] T1027;
  wire[20:0] T5282;
  wire T1028;
  wire T1029;
  wire[20:0] T1030;
  wire[20:0] T1031;
  wire[20:0] T5283;
  wire T1032;
  wire T1033;
  wire[21:0] T1034;
  wire[21:0] T1035;
  wire[21:0] T1036;
  wire[21:0] T5284;
  wire T1037;
  wire T1038;
  wire[21:0] T1039;
  wire[21:0] T1040;
  wire[21:0] T5285;
  wire T1041;
  wire T1042;
  wire[22:0] T1043;
  wire[22:0] T1044;
  wire[22:0] T1045;
  wire[22:0] T5286;
  wire T1046;
  wire T1047;
  wire[22:0] T1048;
  wire[22:0] T1049;
  wire[22:0] T5287;
  wire T1050;
  wire T1051;
  wire[23:0] T1052;
  wire[23:0] T1053;
  wire[23:0] T1054;
  wire[23:0] T5288;
  wire T1055;
  wire T1056;
  wire[23:0] T1057;
  wire[23:0] T1058;
  wire[23:0] T5289;
  wire T1059;
  wire T1060;
  wire[63:0] config_22;
  wire T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire[1:0] G_wire_below_0;
  wire[1:0] G_wire_below_1;
  wire[1:0] G_wire_below_2;
  wire[1:0] G_wire_below_3;
  wire[1:0] H_wire_below_0;
  wire[1:0] H_wire_below_1;
  wire[1:0] H_wire_below_2;
  wire[1:0] H_wire_below_3;
  wire[1:0] H_wire_below_4;
  wire[1:0] H_wire_below_5;
  wire[1:0] H_wire_below_6;
  wire[1:0] H_wire_below_7;
  wire[1:0] H_wire_below_8;
  wire[1:0] H_wire_below_9;
  wire[1:0] H_wire_below_10;
  wire[63:0] config_21;
  wire T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire T1076;
  wire[1:0] H_wire_below_11;
  wire[63:0] config_20;
  wire T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire T1084;
  wire[1:0] H_wire_below_12;
  wire[63:0] config_19;
  wire T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  wire T1090;
  wire T1091;
  wire T1092;
  wire[1:0] H_wire_below_13;
  wire[63:0] config_18;
  wire T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire T1100;
  wire[1:0] H_wire_below_14;
  wire[63:0] config_17;
  wire T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire T1106;
  wire T1107;
  wire T1108;
  wire[1:0] H_wire_below_15;
  wire[63:0] config_16;
  wire T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire T1113;
  wire T1114;
  wire T1115;
  wire T1116;
  wire[1:0] H_wire_below_16;
  wire[63:0] config_15;
  wire T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire T1124;
  wire[1:0] H_wire_below_17;
  wire[63:0] config_14;
  wire T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire T1132;
  wire[1:0] H_wire_below_18;
  wire[63:0] config_13;
  wire T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire[1:0] H_wire_below_19;
  wire[63:0] config_12;
  wire T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire T1145;
  wire T1146;
  wire T1147;
  wire T1148;
  wire[1:0] H_wire_below_20;
  wire[63:0] config_11;
  wire T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire T1153;
  wire T1154;
  wire T1155;
  wire T1156;
  wire[1:0] H_wire_below_21;
  wire[63:0] config_10;
  wire T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire T1164;
  wire[1:0] H_wire_below_22;
  wire[63:0] config_9;
  wire T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire T1169;
  wire T1170;
  wire T1171;
  wire T1172;
  wire[1:0] H_wire_below_23;
  wire[63:0] config_8;
  wire T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire T1180;
  wire[1:0] H_wire_below_24;
  wire[63:0] config_7;
  wire T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire T1185;
  wire T1186;
  wire T1187;
  wire T1188;
  wire[1:0] H_wire_below_25;
  wire[63:0] config_6;
  wire T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire[1:0] H_wire_below_26;
  wire[63:0] config_5;
  wire T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  wire T1204;
  wire[1:0] H_wire_below_27;
  wire[63:0] config_4;
  wire T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire T1209;
  wire T1210;
  wire T1211;
  wire T1212;
  wire[1:0] H_wire_below_28;
  wire[63:0] config_3;
  wire T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire T1217;
  wire T1218;
  wire T1219;
  wire T1220;
  wire[1:0] H_wire_below_29;
  wire[63:0] config_2;
  wire T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  wire T1228;
  wire[1:0] H_wire_below_30;
  wire[63:0] config_1;
  wire T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire T1233;
  wire T1234;
  wire T1235;
  wire T1236;
  wire[1:0] H_wire_below_31;
  wire[63:0] config_0;
  wire T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire[1:0] H_wire_below_32;
  wire[63:0] config_23;
  wire T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire T1257;
  wire T1258;
  wire T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire T1268;
  wire[15:0] V_wire_en_0;
  wire[15:0] T5290;
  wire[16:0] T1269;
  wire[16:0] T1270;
  wire[16:0] T1271;
  wire[16:0] T1272;
  wire[16:0] T1273;
  wire[16:0] T1274;
  wire[16:0] T1275;
  wire[16:0] T1276;
  wire[16:0] T1277;
  wire[16:0] T1278;
  wire[16:0] T1279;
  wire[16:0] T1280;
  wire[16:0] T1281;
  wire[16:0] T1282;
  wire[16:0] T1283;
  wire[16:0] T1284;
  wire[16:0] T1285;
  wire[16:0] T1286;
  wire[16:0] T1287;
  wire[16:0] T5291;
  wire T1288;
  wire T1289;
  wire[16:0] T1290;
  wire[16:0] T1291;
  wire T1292;
  wire T1293;
  wire[3:0] T1294;
  wire T1295;
  wire T1296;
  wire[16:0] T1297;
  wire[16:0] T5292;
  wire[15:0] T1298;
  wire[15:0] T1299;
  wire[15:0] T5293;
  wire T1300;
  wire T1301;
  wire T5294;
  wire[16:0] T1302;
  wire[16:0] T5295;
  wire[15:0] T1303;
  wire T5296;
  wire T1304;
  wire T1305;
  wire[16:0] T1306;
  wire[16:0] T5297;
  wire[14:0] T1307;
  wire[14:0] T1308;
  wire[14:0] T5298;
  wire T1309;
  wire T1310;
  wire[1:0] T5299;
  wire T5300;
  wire[16:0] T1311;
  wire[16:0] T5301;
  wire[14:0] T1312;
  wire[1:0] T5302;
  wire T5303;
  wire T1313;
  wire T1314;
  wire[16:0] T1315;
  wire[16:0] T5304;
  wire[13:0] T1316;
  wire[13:0] T1317;
  wire[13:0] T5305;
  wire T1318;
  wire T1319;
  wire[2:0] T5306;
  wire T5307;
  wire[16:0] T1320;
  wire[16:0] T5308;
  wire[13:0] T1321;
  wire[2:0] T5309;
  wire T5310;
  wire T1322;
  wire T1323;
  wire[16:0] T1324;
  wire[16:0] T5311;
  wire[12:0] T1325;
  wire[12:0] T1326;
  wire[12:0] T5312;
  wire T1327;
  wire T1328;
  wire[3:0] T5313;
  wire T5314;
  wire[16:0] T1329;
  wire[16:0] T5315;
  wire[12:0] T1330;
  wire[3:0] T5316;
  wire T5317;
  wire T1331;
  wire T1332;
  wire[16:0] T1333;
  wire[16:0] T5318;
  wire[11:0] T1334;
  wire[11:0] T1335;
  wire[11:0] T5319;
  wire T1336;
  wire T1337;
  wire[4:0] T5320;
  wire T5321;
  wire[16:0] T1338;
  wire[16:0] T5322;
  wire[11:0] T1339;
  wire[4:0] T5323;
  wire T5324;
  wire T1340;
  wire T1341;
  wire[16:0] T1342;
  wire[16:0] T5325;
  wire[10:0] T1343;
  wire[10:0] T1344;
  wire[10:0] T5326;
  wire T1345;
  wire T1346;
  wire[5:0] T5327;
  wire T5328;
  wire[16:0] T1347;
  wire[16:0] T5329;
  wire[10:0] T1348;
  wire[5:0] T5330;
  wire T5331;
  wire T1349;
  wire T1350;
  wire[16:0] T1351;
  wire[16:0] T5332;
  wire[9:0] T1352;
  wire[9:0] T1353;
  wire[9:0] T5333;
  wire T1354;
  wire T1355;
  wire[6:0] T5334;
  wire T5335;
  wire[16:0] T1356;
  wire[16:0] T5336;
  wire[9:0] T1357;
  wire[6:0] T5337;
  wire T5338;
  wire T1358;
  wire T1359;
  wire[16:0] T1360;
  wire[16:0] T5339;
  wire[8:0] T1361;
  wire[8:0] T1362;
  wire[8:0] T5340;
  wire T1363;
  wire T1364;
  wire[7:0] T5341;
  wire T5342;
  wire[16:0] T1365;
  wire[16:0] T5343;
  wire[8:0] T1366;
  wire[7:0] T5344;
  wire T5345;
  wire T1367;
  wire T1368;
  wire[16:0] T1369;
  wire[16:0] T5346;
  wire[7:0] T1370;
  wire[7:0] T1371;
  wire[7:0] T5347;
  wire T1372;
  wire T1373;
  wire[8:0] T5348;
  wire T5349;
  wire[16:0] T1374;
  wire[16:0] T5350;
  wire[7:0] T1375;
  wire[8:0] T5351;
  wire T5352;
  wire T1376;
  wire T1377;
  wire[16:0] T1378;
  wire[16:0] T5353;
  wire[6:0] T1379;
  wire[6:0] T1380;
  wire[6:0] T5354;
  wire T1381;
  wire T1382;
  wire[9:0] T5355;
  wire T5356;
  wire[16:0] T1383;
  wire[16:0] T5357;
  wire[6:0] T1384;
  wire[9:0] T5358;
  wire T5359;
  wire T1385;
  wire T1386;
  wire[16:0] T1387;
  wire[16:0] T5360;
  wire[5:0] T1388;
  wire[5:0] T1389;
  wire[5:0] T5361;
  wire T1390;
  wire T1391;
  wire[10:0] T5362;
  wire T5363;
  wire[16:0] T1392;
  wire[16:0] T5364;
  wire[5:0] T1393;
  wire[10:0] T5365;
  wire T5366;
  wire T1394;
  wire T1395;
  wire[16:0] T1396;
  wire[16:0] T5367;
  wire[4:0] T1397;
  wire[4:0] T1398;
  wire[4:0] T5368;
  wire T1399;
  wire T1400;
  wire[11:0] T5369;
  wire T5370;
  wire[16:0] T1401;
  wire[16:0] T5371;
  wire[4:0] T1402;
  wire[11:0] T5372;
  wire T5373;
  wire T1403;
  wire T1404;
  wire[16:0] T1405;
  wire[16:0] T5374;
  wire[3:0] T1406;
  wire[3:0] T1407;
  wire[3:0] T5375;
  wire T1408;
  wire T1409;
  wire[12:0] T5376;
  wire T5377;
  wire[16:0] T1410;
  wire[16:0] T5378;
  wire[3:0] T1411;
  wire[12:0] T5379;
  wire T5380;
  wire T1412;
  wire T1413;
  wire[16:0] T1414;
  wire[16:0] T5381;
  wire[2:0] T1415;
  wire[2:0] T1416;
  wire[2:0] T5382;
  wire T1417;
  wire T1418;
  wire[13:0] T5383;
  wire T5384;
  wire[16:0] T1419;
  wire[16:0] T5385;
  wire[2:0] T1420;
  wire[13:0] T5386;
  wire T5387;
  wire T1421;
  wire T1422;
  wire[16:0] T1423;
  wire[16:0] T5388;
  wire[1:0] T1424;
  wire[1:0] T1425;
  wire[1:0] T5389;
  wire T1426;
  wire T1427;
  wire[14:0] T5390;
  wire T5391;
  wire[16:0] T1428;
  wire[16:0] T5392;
  wire[1:0] T1429;
  wire[14:0] T5393;
  wire T5394;
  wire T1430;
  wire T1431;
  wire[15:0] V_wire_en_1;
  wire[15:0] T5395;
  wire[16:0] T1432;
  wire[16:0] T1433;
  wire[16:0] T1434;
  wire[16:0] T1435;
  wire[16:0] T1436;
  wire[16:0] T1437;
  wire[16:0] T1438;
  wire[16:0] T1439;
  wire[16:0] T1440;
  wire[16:0] T1441;
  wire[16:0] T1442;
  wire[16:0] T1443;
  wire[16:0] T1444;
  wire[16:0] T1445;
  wire[16:0] T1446;
  wire[16:0] T1447;
  wire[16:0] T1448;
  wire[16:0] T1449;
  wire[16:0] T1450;
  wire[16:0] T5396;
  wire T1451;
  wire T1452;
  wire[16:0] T1453;
  wire[16:0] T1454;
  wire T1455;
  wire T1456;
  wire[3:0] T1457;
  wire T1458;
  wire T1459;
  wire[16:0] T1460;
  wire[16:0] T5397;
  wire[15:0] T1461;
  wire[15:0] T1462;
  wire[15:0] T5398;
  wire T1463;
  wire T1464;
  wire T5399;
  wire[16:0] T1465;
  wire[16:0] T5400;
  wire[15:0] T1466;
  wire T5401;
  wire T1467;
  wire T1468;
  wire[16:0] T1469;
  wire[16:0] T5402;
  wire[14:0] T1470;
  wire[14:0] T1471;
  wire[14:0] T5403;
  wire T1472;
  wire T1473;
  wire[1:0] T5404;
  wire T5405;
  wire[16:0] T1474;
  wire[16:0] T5406;
  wire[14:0] T1475;
  wire[1:0] T5407;
  wire T5408;
  wire T1476;
  wire T1477;
  wire[16:0] T1478;
  wire[16:0] T5409;
  wire[13:0] T1479;
  wire[13:0] T1480;
  wire[13:0] T5410;
  wire T1481;
  wire T1482;
  wire[2:0] T5411;
  wire T5412;
  wire[16:0] T1483;
  wire[16:0] T5413;
  wire[13:0] T1484;
  wire[2:0] T5414;
  wire T5415;
  wire T1485;
  wire T1486;
  wire[16:0] T1487;
  wire[16:0] T5416;
  wire[12:0] T1488;
  wire[12:0] T1489;
  wire[12:0] T5417;
  wire T1490;
  wire T1491;
  wire[3:0] T5418;
  wire T5419;
  wire[16:0] T1492;
  wire[16:0] T5420;
  wire[12:0] T1493;
  wire[3:0] T5421;
  wire T5422;
  wire T1494;
  wire T1495;
  wire[16:0] T1496;
  wire[16:0] T5423;
  wire[11:0] T1497;
  wire[11:0] T1498;
  wire[11:0] T5424;
  wire T1499;
  wire T1500;
  wire[4:0] T5425;
  wire T5426;
  wire[16:0] T1501;
  wire[16:0] T5427;
  wire[11:0] T1502;
  wire[4:0] T5428;
  wire T5429;
  wire T1503;
  wire T1504;
  wire[16:0] T1505;
  wire[16:0] T5430;
  wire[10:0] T1506;
  wire[10:0] T1507;
  wire[10:0] T5431;
  wire T1508;
  wire T1509;
  wire[5:0] T5432;
  wire T5433;
  wire[16:0] T1510;
  wire[16:0] T5434;
  wire[10:0] T1511;
  wire[5:0] T5435;
  wire T5436;
  wire T1512;
  wire T1513;
  wire[16:0] T1514;
  wire[16:0] T5437;
  wire[9:0] T1515;
  wire[9:0] T1516;
  wire[9:0] T5438;
  wire T1517;
  wire T1518;
  wire[6:0] T5439;
  wire T5440;
  wire[16:0] T1519;
  wire[16:0] T5441;
  wire[9:0] T1520;
  wire[6:0] T5442;
  wire T5443;
  wire T1521;
  wire T1522;
  wire[16:0] T1523;
  wire[16:0] T5444;
  wire[8:0] T1524;
  wire[8:0] T1525;
  wire[8:0] T5445;
  wire T1526;
  wire T1527;
  wire[7:0] T5446;
  wire T5447;
  wire[16:0] T1528;
  wire[16:0] T5448;
  wire[8:0] T1529;
  wire[7:0] T5449;
  wire T5450;
  wire T1530;
  wire T1531;
  wire[16:0] T1532;
  wire[16:0] T5451;
  wire[7:0] T1533;
  wire[7:0] T1534;
  wire[7:0] T5452;
  wire T1535;
  wire T1536;
  wire[8:0] T5453;
  wire T5454;
  wire[16:0] T1537;
  wire[16:0] T5455;
  wire[7:0] T1538;
  wire[8:0] T5456;
  wire T5457;
  wire T1539;
  wire T1540;
  wire[16:0] T1541;
  wire[16:0] T5458;
  wire[6:0] T1542;
  wire[6:0] T1543;
  wire[6:0] T5459;
  wire T1544;
  wire T1545;
  wire[9:0] T5460;
  wire T5461;
  wire[16:0] T1546;
  wire[16:0] T5462;
  wire[6:0] T1547;
  wire[9:0] T5463;
  wire T5464;
  wire T1548;
  wire T1549;
  wire[16:0] T1550;
  wire[16:0] T5465;
  wire[5:0] T1551;
  wire[5:0] T1552;
  wire[5:0] T5466;
  wire T1553;
  wire T1554;
  wire[10:0] T5467;
  wire T5468;
  wire[16:0] T1555;
  wire[16:0] T5469;
  wire[5:0] T1556;
  wire[10:0] T5470;
  wire T5471;
  wire T1557;
  wire T1558;
  wire[16:0] T1559;
  wire[16:0] T5472;
  wire[4:0] T1560;
  wire[4:0] T1561;
  wire[4:0] T5473;
  wire T1562;
  wire T1563;
  wire[11:0] T5474;
  wire T5475;
  wire[16:0] T1564;
  wire[16:0] T5476;
  wire[4:0] T1565;
  wire[11:0] T5477;
  wire T5478;
  wire T1566;
  wire T1567;
  wire[16:0] T1568;
  wire[16:0] T5479;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T5480;
  wire T1571;
  wire T1572;
  wire[12:0] T5481;
  wire T5482;
  wire[16:0] T1573;
  wire[16:0] T5483;
  wire[3:0] T1574;
  wire[12:0] T5484;
  wire T5485;
  wire T1575;
  wire T1576;
  wire[16:0] T1577;
  wire[16:0] T5486;
  wire[2:0] T1578;
  wire[2:0] T1579;
  wire[2:0] T5487;
  wire T1580;
  wire T1581;
  wire[13:0] T5488;
  wire T5489;
  wire[16:0] T1582;
  wire[16:0] T5490;
  wire[2:0] T1583;
  wire[13:0] T5491;
  wire T5492;
  wire T1584;
  wire T1585;
  wire[16:0] T1586;
  wire[16:0] T5493;
  wire[1:0] T1587;
  wire[1:0] T1588;
  wire[1:0] T5494;
  wire T1589;
  wire T1590;
  wire[14:0] T5495;
  wire T5496;
  wire[16:0] T1591;
  wire[16:0] T5497;
  wire[1:0] T1592;
  wire[14:0] T5498;
  wire T5499;
  wire T1593;
  wire T1594;
  wire[15:0] V_wire_en_2;
  wire[15:0] T5500;
  wire[16:0] T1595;
  wire[16:0] T1596;
  wire[16:0] T1597;
  wire[16:0] T1598;
  wire[16:0] T1599;
  wire[16:0] T1600;
  wire[16:0] T1601;
  wire[16:0] T1602;
  wire[16:0] T1603;
  wire[16:0] T1604;
  wire[16:0] T1605;
  wire[16:0] T1606;
  wire[16:0] T1607;
  wire[16:0] T1608;
  wire[16:0] T1609;
  wire[16:0] T1610;
  wire[16:0] T1611;
  wire[16:0] T1612;
  wire[16:0] T1613;
  wire[16:0] T5501;
  wire T1614;
  wire T1615;
  wire[16:0] T1616;
  wire[16:0] T1617;
  wire T1618;
  wire T1619;
  wire[3:0] T1620;
  wire T1621;
  wire T1622;
  wire[16:0] T1623;
  wire[16:0] T5502;
  wire[15:0] T1624;
  wire[15:0] T1625;
  wire[15:0] T5503;
  wire T1626;
  wire T1627;
  wire T5504;
  wire[16:0] T1628;
  wire[16:0] T5505;
  wire[15:0] T1629;
  wire T5506;
  wire T1630;
  wire T1631;
  wire[16:0] T1632;
  wire[16:0] T5507;
  wire[14:0] T1633;
  wire[14:0] T1634;
  wire[14:0] T5508;
  wire T1635;
  wire T1636;
  wire[1:0] T5509;
  wire T5510;
  wire[16:0] T1637;
  wire[16:0] T5511;
  wire[14:0] T1638;
  wire[1:0] T5512;
  wire T5513;
  wire T1639;
  wire T1640;
  wire[16:0] T1641;
  wire[16:0] T5514;
  wire[13:0] T1642;
  wire[13:0] T1643;
  wire[13:0] T5515;
  wire T1644;
  wire T1645;
  wire[2:0] T5516;
  wire T5517;
  wire[16:0] T1646;
  wire[16:0] T5518;
  wire[13:0] T1647;
  wire[2:0] T5519;
  wire T5520;
  wire T1648;
  wire T1649;
  wire[16:0] T1650;
  wire[16:0] T5521;
  wire[12:0] T1651;
  wire[12:0] T1652;
  wire[12:0] T5522;
  wire T1653;
  wire T1654;
  wire[3:0] T5523;
  wire T5524;
  wire[16:0] T1655;
  wire[16:0] T5525;
  wire[12:0] T1656;
  wire[3:0] T5526;
  wire T5527;
  wire T1657;
  wire T1658;
  wire[16:0] T1659;
  wire[16:0] T5528;
  wire[11:0] T1660;
  wire[11:0] T1661;
  wire[11:0] T5529;
  wire T1662;
  wire T1663;
  wire[4:0] T5530;
  wire T5531;
  wire[16:0] T1664;
  wire[16:0] T5532;
  wire[11:0] T1665;
  wire[4:0] T5533;
  wire T5534;
  wire T1666;
  wire T1667;
  wire[16:0] T1668;
  wire[16:0] T5535;
  wire[10:0] T1669;
  wire[10:0] T1670;
  wire[10:0] T5536;
  wire T1671;
  wire T1672;
  wire[5:0] T5537;
  wire T5538;
  wire[16:0] T1673;
  wire[16:0] T5539;
  wire[10:0] T1674;
  wire[5:0] T5540;
  wire T5541;
  wire T1675;
  wire T1676;
  wire[16:0] T1677;
  wire[16:0] T5542;
  wire[9:0] T1678;
  wire[9:0] T1679;
  wire[9:0] T5543;
  wire T1680;
  wire T1681;
  wire[6:0] T5544;
  wire T5545;
  wire[16:0] T1682;
  wire[16:0] T5546;
  wire[9:0] T1683;
  wire[6:0] T5547;
  wire T5548;
  wire T1684;
  wire T1685;
  wire[16:0] T1686;
  wire[16:0] T5549;
  wire[8:0] T1687;
  wire[8:0] T1688;
  wire[8:0] T5550;
  wire T1689;
  wire T1690;
  wire[7:0] T5551;
  wire T5552;
  wire[16:0] T1691;
  wire[16:0] T5553;
  wire[8:0] T1692;
  wire[7:0] T5554;
  wire T5555;
  wire T1693;
  wire T1694;
  wire[16:0] T1695;
  wire[16:0] T5556;
  wire[7:0] T1696;
  wire[7:0] T1697;
  wire[7:0] T5557;
  wire T1698;
  wire T1699;
  wire[8:0] T5558;
  wire T5559;
  wire[16:0] T1700;
  wire[16:0] T5560;
  wire[7:0] T1701;
  wire[8:0] T5561;
  wire T5562;
  wire T1702;
  wire T1703;
  wire[16:0] T1704;
  wire[16:0] T5563;
  wire[6:0] T1705;
  wire[6:0] T1706;
  wire[6:0] T5564;
  wire T1707;
  wire T1708;
  wire[9:0] T5565;
  wire T5566;
  wire[16:0] T1709;
  wire[16:0] T5567;
  wire[6:0] T1710;
  wire[9:0] T5568;
  wire T5569;
  wire T1711;
  wire T1712;
  wire[16:0] T1713;
  wire[16:0] T5570;
  wire[5:0] T1714;
  wire[5:0] T1715;
  wire[5:0] T5571;
  wire T1716;
  wire T1717;
  wire[10:0] T5572;
  wire T5573;
  wire[16:0] T1718;
  wire[16:0] T5574;
  wire[5:0] T1719;
  wire[10:0] T5575;
  wire T5576;
  wire T1720;
  wire T1721;
  wire[16:0] T1722;
  wire[16:0] T5577;
  wire[4:0] T1723;
  wire[4:0] T1724;
  wire[4:0] T5578;
  wire T1725;
  wire T1726;
  wire[11:0] T5579;
  wire T5580;
  wire[16:0] T1727;
  wire[16:0] T5581;
  wire[4:0] T1728;
  wire[11:0] T5582;
  wire T5583;
  wire T1729;
  wire T1730;
  wire[16:0] T1731;
  wire[16:0] T5584;
  wire[3:0] T1732;
  wire[3:0] T1733;
  wire[3:0] T5585;
  wire T1734;
  wire T1735;
  wire[12:0] T5586;
  wire T5587;
  wire[16:0] T1736;
  wire[16:0] T5588;
  wire[3:0] T1737;
  wire[12:0] T5589;
  wire T5590;
  wire T1738;
  wire T1739;
  wire[16:0] T1740;
  wire[16:0] T5591;
  wire[2:0] T1741;
  wire[2:0] T1742;
  wire[2:0] T5592;
  wire T1743;
  wire T1744;
  wire[13:0] T5593;
  wire T5594;
  wire[16:0] T1745;
  wire[16:0] T5595;
  wire[2:0] T1746;
  wire[13:0] T5596;
  wire T5597;
  wire T1747;
  wire T1748;
  wire[16:0] T1749;
  wire[16:0] T5598;
  wire[1:0] T1750;
  wire[1:0] T1751;
  wire[1:0] T5599;
  wire T1752;
  wire T1753;
  wire[14:0] T5600;
  wire T5601;
  wire[16:0] T1754;
  wire[16:0] T5602;
  wire[1:0] T1755;
  wire[14:0] T5603;
  wire T5604;
  wire T1756;
  wire T1757;
  wire[15:0] V_wire_en_3;
  wire[15:0] T5605;
  wire[16:0] T1758;
  wire[16:0] T1759;
  wire[16:0] T1760;
  wire[16:0] T1761;
  wire[16:0] T1762;
  wire[16:0] T1763;
  wire[16:0] T1764;
  wire[16:0] T1765;
  wire[16:0] T1766;
  wire[16:0] T1767;
  wire[16:0] T1768;
  wire[16:0] T1769;
  wire[16:0] T1770;
  wire[16:0] T1771;
  wire[16:0] T1772;
  wire[16:0] T1773;
  wire[16:0] T1774;
  wire[16:0] T1775;
  wire[16:0] T1776;
  wire[16:0] T5606;
  wire T1777;
  wire T1778;
  wire[16:0] T1779;
  wire[16:0] T1780;
  wire T1781;
  wire T1782;
  wire[3:0] T1783;
  wire T1784;
  wire T1785;
  wire[16:0] T1786;
  wire[16:0] T5607;
  wire[15:0] T1787;
  wire[15:0] T1788;
  wire[15:0] T5608;
  wire T1789;
  wire T1790;
  wire T5609;
  wire[16:0] T1791;
  wire[16:0] T5610;
  wire[15:0] T1792;
  wire T5611;
  wire T1793;
  wire T1794;
  wire[16:0] T1795;
  wire[16:0] T5612;
  wire[14:0] T1796;
  wire[14:0] T1797;
  wire[14:0] T5613;
  wire T1798;
  wire T1799;
  wire[1:0] T5614;
  wire T5615;
  wire[16:0] T1800;
  wire[16:0] T5616;
  wire[14:0] T1801;
  wire[1:0] T5617;
  wire T5618;
  wire T1802;
  wire T1803;
  wire[16:0] T1804;
  wire[16:0] T5619;
  wire[13:0] T1805;
  wire[13:0] T1806;
  wire[13:0] T5620;
  wire T1807;
  wire T1808;
  wire[2:0] T5621;
  wire T5622;
  wire[16:0] T1809;
  wire[16:0] T5623;
  wire[13:0] T1810;
  wire[2:0] T5624;
  wire T5625;
  wire T1811;
  wire T1812;
  wire[16:0] T1813;
  wire[16:0] T5626;
  wire[12:0] T1814;
  wire[12:0] T1815;
  wire[12:0] T5627;
  wire T1816;
  wire T1817;
  wire[3:0] T5628;
  wire T5629;
  wire[16:0] T1818;
  wire[16:0] T5630;
  wire[12:0] T1819;
  wire[3:0] T5631;
  wire T5632;
  wire T1820;
  wire T1821;
  wire[16:0] T1822;
  wire[16:0] T5633;
  wire[11:0] T1823;
  wire[11:0] T1824;
  wire[11:0] T5634;
  wire T1825;
  wire T1826;
  wire[4:0] T5635;
  wire T5636;
  wire[16:0] T1827;
  wire[16:0] T5637;
  wire[11:0] T1828;
  wire[4:0] T5638;
  wire T5639;
  wire T1829;
  wire T1830;
  wire[16:0] T1831;
  wire[16:0] T5640;
  wire[10:0] T1832;
  wire[10:0] T1833;
  wire[10:0] T5641;
  wire T1834;
  wire T1835;
  wire[5:0] T5642;
  wire T5643;
  wire[16:0] T1836;
  wire[16:0] T5644;
  wire[10:0] T1837;
  wire[5:0] T5645;
  wire T5646;
  wire T1838;
  wire T1839;
  wire[16:0] T1840;
  wire[16:0] T5647;
  wire[9:0] T1841;
  wire[9:0] T1842;
  wire[9:0] T5648;
  wire T1843;
  wire T1844;
  wire[6:0] T5649;
  wire T5650;
  wire[16:0] T1845;
  wire[16:0] T5651;
  wire[9:0] T1846;
  wire[6:0] T5652;
  wire T5653;
  wire T1847;
  wire T1848;
  wire[16:0] T1849;
  wire[16:0] T5654;
  wire[8:0] T1850;
  wire[8:0] T1851;
  wire[8:0] T5655;
  wire T1852;
  wire T1853;
  wire[7:0] T5656;
  wire T5657;
  wire[16:0] T1854;
  wire[16:0] T5658;
  wire[8:0] T1855;
  wire[7:0] T5659;
  wire T5660;
  wire T1856;
  wire T1857;
  wire[16:0] T1858;
  wire[16:0] T5661;
  wire[7:0] T1859;
  wire[7:0] T1860;
  wire[7:0] T5662;
  wire T1861;
  wire T1862;
  wire[8:0] T5663;
  wire T5664;
  wire[16:0] T1863;
  wire[16:0] T5665;
  wire[7:0] T1864;
  wire[8:0] T5666;
  wire T5667;
  wire T1865;
  wire T1866;
  wire[16:0] T1867;
  wire[16:0] T5668;
  wire[6:0] T1868;
  wire[6:0] T1869;
  wire[6:0] T5669;
  wire T1870;
  wire T1871;
  wire[9:0] T5670;
  wire T5671;
  wire[16:0] T1872;
  wire[16:0] T5672;
  wire[6:0] T1873;
  wire[9:0] T5673;
  wire T5674;
  wire T1874;
  wire T1875;
  wire[16:0] T1876;
  wire[16:0] T5675;
  wire[5:0] T1877;
  wire[5:0] T1878;
  wire[5:0] T5676;
  wire T1879;
  wire T1880;
  wire[10:0] T5677;
  wire T5678;
  wire[16:0] T1881;
  wire[16:0] T5679;
  wire[5:0] T1882;
  wire[10:0] T5680;
  wire T5681;
  wire T1883;
  wire T1884;
  wire[16:0] T1885;
  wire[16:0] T5682;
  wire[4:0] T1886;
  wire[4:0] T1887;
  wire[4:0] T5683;
  wire T1888;
  wire T1889;
  wire[11:0] T5684;
  wire T5685;
  wire[16:0] T1890;
  wire[16:0] T5686;
  wire[4:0] T1891;
  wire[11:0] T5687;
  wire T5688;
  wire T1892;
  wire T1893;
  wire[16:0] T1894;
  wire[16:0] T5689;
  wire[3:0] T1895;
  wire[3:0] T1896;
  wire[3:0] T5690;
  wire T1897;
  wire T1898;
  wire[12:0] T5691;
  wire T5692;
  wire[16:0] T1899;
  wire[16:0] T5693;
  wire[3:0] T1900;
  wire[12:0] T5694;
  wire T5695;
  wire T1901;
  wire T1902;
  wire[16:0] T1903;
  wire[16:0] T5696;
  wire[2:0] T1904;
  wire[2:0] T1905;
  wire[2:0] T5697;
  wire T1906;
  wire T1907;
  wire[13:0] T5698;
  wire T5699;
  wire[16:0] T1908;
  wire[16:0] T5700;
  wire[2:0] T1909;
  wire[13:0] T5701;
  wire T5702;
  wire T1910;
  wire T1911;
  wire[16:0] T1912;
  wire[16:0] T5703;
  wire[1:0] T1913;
  wire[1:0] T1914;
  wire[1:0] T5704;
  wire T1915;
  wire T1916;
  wire[14:0] T5705;
  wire T5706;
  wire[16:0] T1917;
  wire[16:0] T5707;
  wire[1:0] T1918;
  wire[14:0] T5708;
  wire T5709;
  wire T1919;
  wire T1920;
  wire[15:0] V_wire_en_4;
  wire[15:0] T5710;
  wire[16:0] T1921;
  wire[16:0] T1922;
  wire[16:0] T1923;
  wire[16:0] T1924;
  wire[16:0] T1925;
  wire[16:0] T1926;
  wire[16:0] T1927;
  wire[16:0] T1928;
  wire[16:0] T1929;
  wire[16:0] T1930;
  wire[16:0] T1931;
  wire[16:0] T1932;
  wire[16:0] T1933;
  wire[16:0] T1934;
  wire[16:0] T1935;
  wire[16:0] T1936;
  wire[16:0] T1937;
  wire[16:0] T1938;
  wire[16:0] T1939;
  wire[16:0] T5711;
  wire T1940;
  wire T1941;
  wire[16:0] T1942;
  wire[16:0] T1943;
  wire T1944;
  wire T1945;
  wire[3:0] T1946;
  wire T1947;
  wire T1948;
  wire[16:0] T1949;
  wire[16:0] T5712;
  wire[15:0] T1950;
  wire[15:0] T1951;
  wire[15:0] T5713;
  wire T1952;
  wire T1953;
  wire T5714;
  wire[16:0] T1954;
  wire[16:0] T5715;
  wire[15:0] T1955;
  wire T5716;
  wire T1956;
  wire T1957;
  wire[16:0] T1958;
  wire[16:0] T5717;
  wire[14:0] T1959;
  wire[14:0] T1960;
  wire[14:0] T5718;
  wire T1961;
  wire T1962;
  wire[1:0] T5719;
  wire T5720;
  wire[16:0] T1963;
  wire[16:0] T5721;
  wire[14:0] T1964;
  wire[1:0] T5722;
  wire T5723;
  wire T1965;
  wire T1966;
  wire[16:0] T1967;
  wire[16:0] T5724;
  wire[13:0] T1968;
  wire[13:0] T1969;
  wire[13:0] T5725;
  wire T1970;
  wire T1971;
  wire[2:0] T5726;
  wire T5727;
  wire[16:0] T1972;
  wire[16:0] T5728;
  wire[13:0] T1973;
  wire[2:0] T5729;
  wire T5730;
  wire T1974;
  wire T1975;
  wire[16:0] T1976;
  wire[16:0] T5731;
  wire[12:0] T1977;
  wire[12:0] T1978;
  wire[12:0] T5732;
  wire T1979;
  wire T1980;
  wire[3:0] T5733;
  wire T5734;
  wire[16:0] T1981;
  wire[16:0] T5735;
  wire[12:0] T1982;
  wire[3:0] T5736;
  wire T5737;
  wire T1983;
  wire T1984;
  wire[16:0] T1985;
  wire[16:0] T5738;
  wire[11:0] T1986;
  wire[11:0] T1987;
  wire[11:0] T5739;
  wire T1988;
  wire T1989;
  wire[4:0] T5740;
  wire T5741;
  wire[16:0] T1990;
  wire[16:0] T5742;
  wire[11:0] T1991;
  wire[4:0] T5743;
  wire T5744;
  wire T1992;
  wire T1993;
  wire[16:0] T1994;
  wire[16:0] T5745;
  wire[10:0] T1995;
  wire[10:0] T1996;
  wire[10:0] T5746;
  wire T1997;
  wire T1998;
  wire[5:0] T5747;
  wire T5748;
  wire[16:0] T1999;
  wire[16:0] T5749;
  wire[10:0] T2000;
  wire[5:0] T5750;
  wire T5751;
  wire T2001;
  wire T2002;
  wire[16:0] T2003;
  wire[16:0] T5752;
  wire[9:0] T2004;
  wire[9:0] T2005;
  wire[9:0] T5753;
  wire T2006;
  wire T2007;
  wire[6:0] T5754;
  wire T5755;
  wire[16:0] T2008;
  wire[16:0] T5756;
  wire[9:0] T2009;
  wire[6:0] T5757;
  wire T5758;
  wire T2010;
  wire T2011;
  wire[16:0] T2012;
  wire[16:0] T5759;
  wire[8:0] T2013;
  wire[8:0] T2014;
  wire[8:0] T5760;
  wire T2015;
  wire T2016;
  wire[7:0] T5761;
  wire T5762;
  wire[16:0] T2017;
  wire[16:0] T5763;
  wire[8:0] T2018;
  wire[7:0] T5764;
  wire T5765;
  wire T2019;
  wire T2020;
  wire[16:0] T2021;
  wire[16:0] T5766;
  wire[7:0] T2022;
  wire[7:0] T2023;
  wire[7:0] T5767;
  wire T2024;
  wire T2025;
  wire[8:0] T5768;
  wire T5769;
  wire[16:0] T2026;
  wire[16:0] T5770;
  wire[7:0] T2027;
  wire[8:0] T5771;
  wire T5772;
  wire T2028;
  wire T2029;
  wire[16:0] T2030;
  wire[16:0] T5773;
  wire[6:0] T2031;
  wire[6:0] T2032;
  wire[6:0] T5774;
  wire T2033;
  wire T2034;
  wire[9:0] T5775;
  wire T5776;
  wire[16:0] T2035;
  wire[16:0] T5777;
  wire[6:0] T2036;
  wire[9:0] T5778;
  wire T5779;
  wire T2037;
  wire T2038;
  wire[16:0] T2039;
  wire[16:0] T5780;
  wire[5:0] T2040;
  wire[5:0] T2041;
  wire[5:0] T5781;
  wire T2042;
  wire T2043;
  wire[10:0] T5782;
  wire T5783;
  wire[16:0] T2044;
  wire[16:0] T5784;
  wire[5:0] T2045;
  wire[10:0] T5785;
  wire T5786;
  wire T2046;
  wire T2047;
  wire[16:0] T2048;
  wire[16:0] T5787;
  wire[4:0] T2049;
  wire[4:0] T2050;
  wire[4:0] T5788;
  wire T2051;
  wire T2052;
  wire[11:0] T5789;
  wire T5790;
  wire[16:0] T2053;
  wire[16:0] T5791;
  wire[4:0] T2054;
  wire[11:0] T5792;
  wire T5793;
  wire T2055;
  wire T2056;
  wire[16:0] T2057;
  wire[16:0] T5794;
  wire[3:0] T2058;
  wire[3:0] T2059;
  wire[3:0] T5795;
  wire T2060;
  wire T2061;
  wire[12:0] T5796;
  wire T5797;
  wire[16:0] T2062;
  wire[16:0] T5798;
  wire[3:0] T2063;
  wire[12:0] T5799;
  wire T5800;
  wire T2064;
  wire T2065;
  wire[16:0] T2066;
  wire[16:0] T5801;
  wire[2:0] T2067;
  wire[2:0] T2068;
  wire[2:0] T5802;
  wire T2069;
  wire T2070;
  wire[13:0] T5803;
  wire T5804;
  wire[16:0] T2071;
  wire[16:0] T5805;
  wire[2:0] T2072;
  wire[13:0] T5806;
  wire T5807;
  wire T2073;
  wire T2074;
  wire[16:0] T2075;
  wire[16:0] T5808;
  wire[1:0] T2076;
  wire[1:0] T2077;
  wire[1:0] T5809;
  wire T2078;
  wire T2079;
  wire[14:0] T5810;
  wire T5811;
  wire[16:0] T2080;
  wire[16:0] T5812;
  wire[1:0] T2081;
  wire[14:0] T5813;
  wire T5814;
  wire T2082;
  wire T2083;
  wire[15:0] V_wire_en_5;
  wire[15:0] T5815;
  wire[16:0] T2084;
  wire[16:0] T2085;
  wire[16:0] T2086;
  wire[16:0] T2087;
  wire[16:0] T2088;
  wire[16:0] T2089;
  wire[16:0] T2090;
  wire[16:0] T2091;
  wire[16:0] T2092;
  wire[16:0] T2093;
  wire[16:0] T2094;
  wire[16:0] T2095;
  wire[16:0] T2096;
  wire[16:0] T2097;
  wire[16:0] T2098;
  wire[16:0] T2099;
  wire[16:0] T2100;
  wire[16:0] T2101;
  wire[16:0] T2102;
  wire[16:0] T5816;
  wire T2103;
  wire T2104;
  wire[16:0] T2105;
  wire[16:0] T2106;
  wire T2107;
  wire T2108;
  wire[3:0] T2109;
  wire T2110;
  wire T2111;
  wire[16:0] T2112;
  wire[16:0] T5817;
  wire[15:0] T2113;
  wire[15:0] T2114;
  wire[15:0] T5818;
  wire T2115;
  wire T2116;
  wire T5819;
  wire[16:0] T2117;
  wire[16:0] T5820;
  wire[15:0] T2118;
  wire T5821;
  wire T2119;
  wire T2120;
  wire[16:0] T2121;
  wire[16:0] T5822;
  wire[14:0] T2122;
  wire[14:0] T2123;
  wire[14:0] T5823;
  wire T2124;
  wire T2125;
  wire[1:0] T5824;
  wire T5825;
  wire[16:0] T2126;
  wire[16:0] T5826;
  wire[14:0] T2127;
  wire[1:0] T5827;
  wire T5828;
  wire T2128;
  wire T2129;
  wire[16:0] T2130;
  wire[16:0] T5829;
  wire[13:0] T2131;
  wire[13:0] T2132;
  wire[13:0] T5830;
  wire T2133;
  wire T2134;
  wire[2:0] T5831;
  wire T5832;
  wire[16:0] T2135;
  wire[16:0] T5833;
  wire[13:0] T2136;
  wire[2:0] T5834;
  wire T5835;
  wire T2137;
  wire T2138;
  wire[16:0] T2139;
  wire[16:0] T5836;
  wire[12:0] T2140;
  wire[12:0] T2141;
  wire[12:0] T5837;
  wire T2142;
  wire T2143;
  wire[3:0] T5838;
  wire T5839;
  wire[16:0] T2144;
  wire[16:0] T5840;
  wire[12:0] T2145;
  wire[3:0] T5841;
  wire T5842;
  wire T2146;
  wire T2147;
  wire[16:0] T2148;
  wire[16:0] T5843;
  wire[11:0] T2149;
  wire[11:0] T2150;
  wire[11:0] T5844;
  wire T2151;
  wire T2152;
  wire[4:0] T5845;
  wire T5846;
  wire[16:0] T2153;
  wire[16:0] T5847;
  wire[11:0] T2154;
  wire[4:0] T5848;
  wire T5849;
  wire T2155;
  wire T2156;
  wire[16:0] T2157;
  wire[16:0] T5850;
  wire[10:0] T2158;
  wire[10:0] T2159;
  wire[10:0] T5851;
  wire T2160;
  wire T2161;
  wire[5:0] T5852;
  wire T5853;
  wire[16:0] T2162;
  wire[16:0] T5854;
  wire[10:0] T2163;
  wire[5:0] T5855;
  wire T5856;
  wire T2164;
  wire T2165;
  wire[16:0] T2166;
  wire[16:0] T5857;
  wire[9:0] T2167;
  wire[9:0] T2168;
  wire[9:0] T5858;
  wire T2169;
  wire T2170;
  wire[6:0] T5859;
  wire T5860;
  wire[16:0] T2171;
  wire[16:0] T5861;
  wire[9:0] T2172;
  wire[6:0] T5862;
  wire T5863;
  wire T2173;
  wire T2174;
  wire[16:0] T2175;
  wire[16:0] T5864;
  wire[8:0] T2176;
  wire[8:0] T2177;
  wire[8:0] T5865;
  wire T2178;
  wire T2179;
  wire[7:0] T5866;
  wire T5867;
  wire[16:0] T2180;
  wire[16:0] T5868;
  wire[8:0] T2181;
  wire[7:0] T5869;
  wire T5870;
  wire T2182;
  wire T2183;
  wire[16:0] T2184;
  wire[16:0] T5871;
  wire[7:0] T2185;
  wire[7:0] T2186;
  wire[7:0] T5872;
  wire T2187;
  wire T2188;
  wire[8:0] T5873;
  wire T5874;
  wire[16:0] T2189;
  wire[16:0] T5875;
  wire[7:0] T2190;
  wire[8:0] T5876;
  wire T5877;
  wire T2191;
  wire T2192;
  wire[16:0] T2193;
  wire[16:0] T5878;
  wire[6:0] T2194;
  wire[6:0] T2195;
  wire[6:0] T5879;
  wire T2196;
  wire T2197;
  wire[9:0] T5880;
  wire T5881;
  wire[16:0] T2198;
  wire[16:0] T5882;
  wire[6:0] T2199;
  wire[9:0] T5883;
  wire T5884;
  wire T2200;
  wire T2201;
  wire[16:0] T2202;
  wire[16:0] T5885;
  wire[5:0] T2203;
  wire[5:0] T2204;
  wire[5:0] T5886;
  wire T2205;
  wire T2206;
  wire[10:0] T5887;
  wire T5888;
  wire[16:0] T2207;
  wire[16:0] T5889;
  wire[5:0] T2208;
  wire[10:0] T5890;
  wire T5891;
  wire T2209;
  wire T2210;
  wire[16:0] T2211;
  wire[16:0] T5892;
  wire[4:0] T2212;
  wire[4:0] T2213;
  wire[4:0] T5893;
  wire T2214;
  wire T2215;
  wire[11:0] T5894;
  wire T5895;
  wire[16:0] T2216;
  wire[16:0] T5896;
  wire[4:0] T2217;
  wire[11:0] T5897;
  wire T5898;
  wire T2218;
  wire T2219;
  wire[16:0] T2220;
  wire[16:0] T5899;
  wire[3:0] T2221;
  wire[3:0] T2222;
  wire[3:0] T5900;
  wire T2223;
  wire T2224;
  wire[12:0] T5901;
  wire T5902;
  wire[16:0] T2225;
  wire[16:0] T5903;
  wire[3:0] T2226;
  wire[12:0] T5904;
  wire T5905;
  wire T2227;
  wire T2228;
  wire[16:0] T2229;
  wire[16:0] T5906;
  wire[2:0] T2230;
  wire[2:0] T2231;
  wire[2:0] T5907;
  wire T2232;
  wire T2233;
  wire[13:0] T5908;
  wire T5909;
  wire[16:0] T2234;
  wire[16:0] T5910;
  wire[2:0] T2235;
  wire[13:0] T5911;
  wire T5912;
  wire T2236;
  wire T2237;
  wire[16:0] T2238;
  wire[16:0] T5913;
  wire[1:0] T2239;
  wire[1:0] T2240;
  wire[1:0] T5914;
  wire T2241;
  wire T2242;
  wire[14:0] T5915;
  wire T5916;
  wire[16:0] T2243;
  wire[16:0] T5917;
  wire[1:0] T2244;
  wire[14:0] T5918;
  wire T5919;
  wire T2245;
  wire T2246;
  wire[15:0] V_wire_en_6;
  wire[15:0] T5920;
  wire[16:0] T2247;
  wire[16:0] T2248;
  wire[16:0] T2249;
  wire[16:0] T2250;
  wire[16:0] T2251;
  wire[16:0] T2252;
  wire[16:0] T2253;
  wire[16:0] T2254;
  wire[16:0] T2255;
  wire[16:0] T2256;
  wire[16:0] T2257;
  wire[16:0] T2258;
  wire[16:0] T2259;
  wire[16:0] T2260;
  wire[16:0] T2261;
  wire[16:0] T2262;
  wire[16:0] T2263;
  wire[16:0] T2264;
  wire[16:0] T2265;
  wire[16:0] T5921;
  wire T2266;
  wire T2267;
  wire[16:0] T2268;
  wire[16:0] T2269;
  wire T2270;
  wire T2271;
  wire[3:0] T2272;
  wire T2273;
  wire T2274;
  wire[16:0] T2275;
  wire[16:0] T5922;
  wire[15:0] T2276;
  wire[15:0] T2277;
  wire[15:0] T5923;
  wire T2278;
  wire T2279;
  wire T5924;
  wire[16:0] T2280;
  wire[16:0] T5925;
  wire[15:0] T2281;
  wire T5926;
  wire T2282;
  wire T2283;
  wire[16:0] T2284;
  wire[16:0] T5927;
  wire[14:0] T2285;
  wire[14:0] T2286;
  wire[14:0] T5928;
  wire T2287;
  wire T2288;
  wire[1:0] T5929;
  wire T5930;
  wire[16:0] T2289;
  wire[16:0] T5931;
  wire[14:0] T2290;
  wire[1:0] T5932;
  wire T5933;
  wire T2291;
  wire T2292;
  wire[16:0] T2293;
  wire[16:0] T5934;
  wire[13:0] T2294;
  wire[13:0] T2295;
  wire[13:0] T5935;
  wire T2296;
  wire T2297;
  wire[2:0] T5936;
  wire T5937;
  wire[16:0] T2298;
  wire[16:0] T5938;
  wire[13:0] T2299;
  wire[2:0] T5939;
  wire T5940;
  wire T2300;
  wire T2301;
  wire[16:0] T2302;
  wire[16:0] T5941;
  wire[12:0] T2303;
  wire[12:0] T2304;
  wire[12:0] T5942;
  wire T2305;
  wire T2306;
  wire[3:0] T5943;
  wire T5944;
  wire[16:0] T2307;
  wire[16:0] T5945;
  wire[12:0] T2308;
  wire[3:0] T5946;
  wire T5947;
  wire T2309;
  wire T2310;
  wire[16:0] T2311;
  wire[16:0] T5948;
  wire[11:0] T2312;
  wire[11:0] T2313;
  wire[11:0] T5949;
  wire T2314;
  wire T2315;
  wire[4:0] T5950;
  wire T5951;
  wire[16:0] T2316;
  wire[16:0] T5952;
  wire[11:0] T2317;
  wire[4:0] T5953;
  wire T5954;
  wire T2318;
  wire T2319;
  wire[16:0] T2320;
  wire[16:0] T5955;
  wire[10:0] T2321;
  wire[10:0] T2322;
  wire[10:0] T5956;
  wire T2323;
  wire T2324;
  wire[5:0] T5957;
  wire T5958;
  wire[16:0] T2325;
  wire[16:0] T5959;
  wire[10:0] T2326;
  wire[5:0] T5960;
  wire T5961;
  wire T2327;
  wire T2328;
  wire[16:0] T2329;
  wire[16:0] T5962;
  wire[9:0] T2330;
  wire[9:0] T2331;
  wire[9:0] T5963;
  wire T2332;
  wire T2333;
  wire[6:0] T5964;
  wire T5965;
  wire[16:0] T2334;
  wire[16:0] T5966;
  wire[9:0] T2335;
  wire[6:0] T5967;
  wire T5968;
  wire T2336;
  wire T2337;
  wire[16:0] T2338;
  wire[16:0] T5969;
  wire[8:0] T2339;
  wire[8:0] T2340;
  wire[8:0] T5970;
  wire T2341;
  wire T2342;
  wire[7:0] T5971;
  wire T5972;
  wire[16:0] T2343;
  wire[16:0] T5973;
  wire[8:0] T2344;
  wire[7:0] T5974;
  wire T5975;
  wire T2345;
  wire T2346;
  wire[16:0] T2347;
  wire[16:0] T5976;
  wire[7:0] T2348;
  wire[7:0] T2349;
  wire[7:0] T5977;
  wire T2350;
  wire T2351;
  wire[8:0] T5978;
  wire T5979;
  wire[16:0] T2352;
  wire[16:0] T5980;
  wire[7:0] T2353;
  wire[8:0] T5981;
  wire T5982;
  wire T2354;
  wire T2355;
  wire[16:0] T2356;
  wire[16:0] T5983;
  wire[6:0] T2357;
  wire[6:0] T2358;
  wire[6:0] T5984;
  wire T2359;
  wire T2360;
  wire[9:0] T5985;
  wire T5986;
  wire[16:0] T2361;
  wire[16:0] T5987;
  wire[6:0] T2362;
  wire[9:0] T5988;
  wire T5989;
  wire T2363;
  wire T2364;
  wire[16:0] T2365;
  wire[16:0] T5990;
  wire[5:0] T2366;
  wire[5:0] T2367;
  wire[5:0] T5991;
  wire T2368;
  wire T2369;
  wire[10:0] T5992;
  wire T5993;
  wire[16:0] T2370;
  wire[16:0] T5994;
  wire[5:0] T2371;
  wire[10:0] T5995;
  wire T5996;
  wire T2372;
  wire T2373;
  wire[16:0] T2374;
  wire[16:0] T5997;
  wire[4:0] T2375;
  wire[4:0] T2376;
  wire[4:0] T5998;
  wire T2377;
  wire T2378;
  wire[11:0] T5999;
  wire T6000;
  wire[16:0] T2379;
  wire[16:0] T6001;
  wire[4:0] T2380;
  wire[11:0] T6002;
  wire T6003;
  wire T2381;
  wire T2382;
  wire[16:0] T2383;
  wire[16:0] T6004;
  wire[3:0] T2384;
  wire[3:0] T2385;
  wire[3:0] T6005;
  wire T2386;
  wire T2387;
  wire[12:0] T6006;
  wire T6007;
  wire[16:0] T2388;
  wire[16:0] T6008;
  wire[3:0] T2389;
  wire[12:0] T6009;
  wire T6010;
  wire T2390;
  wire T2391;
  wire[16:0] T2392;
  wire[16:0] T6011;
  wire[2:0] T2393;
  wire[2:0] T2394;
  wire[2:0] T6012;
  wire T2395;
  wire T2396;
  wire[13:0] T6013;
  wire T6014;
  wire[16:0] T2397;
  wire[16:0] T6015;
  wire[2:0] T2398;
  wire[13:0] T6016;
  wire T6017;
  wire T2399;
  wire T2400;
  wire[16:0] T2401;
  wire[16:0] T6018;
  wire[1:0] T2402;
  wire[1:0] T2403;
  wire[1:0] T6019;
  wire T2404;
  wire T2405;
  wire[14:0] T6020;
  wire T6021;
  wire[16:0] T2406;
  wire[16:0] T6022;
  wire[1:0] T2407;
  wire[14:0] T6023;
  wire T6024;
  wire T2408;
  wire T2409;
  wire[15:0] V_wire_en_7;
  wire[15:0] T6025;
  wire[16:0] T2410;
  wire[16:0] T2411;
  wire[16:0] T2412;
  wire[16:0] T2413;
  wire[16:0] T2414;
  wire[16:0] T2415;
  wire[16:0] T2416;
  wire[16:0] T2417;
  wire[16:0] T2418;
  wire[16:0] T2419;
  wire[16:0] T2420;
  wire[16:0] T2421;
  wire[16:0] T2422;
  wire[16:0] T2423;
  wire[16:0] T2424;
  wire[16:0] T2425;
  wire[16:0] T2426;
  wire[16:0] T2427;
  wire[16:0] T2428;
  wire[16:0] T6026;
  wire T2429;
  wire T2430;
  wire[16:0] T2431;
  wire[16:0] T2432;
  wire T2433;
  wire T2434;
  wire[3:0] T2435;
  wire T2436;
  wire T2437;
  wire[16:0] T2438;
  wire[16:0] T6027;
  wire[15:0] T2439;
  wire[15:0] T2440;
  wire[15:0] T6028;
  wire T2441;
  wire T2442;
  wire T6029;
  wire[16:0] T2443;
  wire[16:0] T6030;
  wire[15:0] T2444;
  wire T6031;
  wire T2445;
  wire T2446;
  wire[16:0] T2447;
  wire[16:0] T6032;
  wire[14:0] T2448;
  wire[14:0] T2449;
  wire[14:0] T6033;
  wire T2450;
  wire T2451;
  wire[1:0] T6034;
  wire T6035;
  wire[16:0] T2452;
  wire[16:0] T6036;
  wire[14:0] T2453;
  wire[1:0] T6037;
  wire T6038;
  wire T2454;
  wire T2455;
  wire[16:0] T2456;
  wire[16:0] T6039;
  wire[13:0] T2457;
  wire[13:0] T2458;
  wire[13:0] T6040;
  wire T2459;
  wire T2460;
  wire[2:0] T6041;
  wire T6042;
  wire[16:0] T2461;
  wire[16:0] T6043;
  wire[13:0] T2462;
  wire[2:0] T6044;
  wire T6045;
  wire T2463;
  wire T2464;
  wire[16:0] T2465;
  wire[16:0] T6046;
  wire[12:0] T2466;
  wire[12:0] T2467;
  wire[12:0] T6047;
  wire T2468;
  wire T2469;
  wire[3:0] T6048;
  wire T6049;
  wire[16:0] T2470;
  wire[16:0] T6050;
  wire[12:0] T2471;
  wire[3:0] T6051;
  wire T6052;
  wire T2472;
  wire T2473;
  wire[16:0] T2474;
  wire[16:0] T6053;
  wire[11:0] T2475;
  wire[11:0] T2476;
  wire[11:0] T6054;
  wire T2477;
  wire T2478;
  wire[4:0] T6055;
  wire T6056;
  wire[16:0] T2479;
  wire[16:0] T6057;
  wire[11:0] T2480;
  wire[4:0] T6058;
  wire T6059;
  wire T2481;
  wire T2482;
  wire[16:0] T2483;
  wire[16:0] T6060;
  wire[10:0] T2484;
  wire[10:0] T2485;
  wire[10:0] T6061;
  wire T2486;
  wire T2487;
  wire[5:0] T6062;
  wire T6063;
  wire[16:0] T2488;
  wire[16:0] T6064;
  wire[10:0] T2489;
  wire[5:0] T6065;
  wire T6066;
  wire T2490;
  wire T2491;
  wire[16:0] T2492;
  wire[16:0] T6067;
  wire[9:0] T2493;
  wire[9:0] T2494;
  wire[9:0] T6068;
  wire T2495;
  wire T2496;
  wire[6:0] T6069;
  wire T6070;
  wire[16:0] T2497;
  wire[16:0] T6071;
  wire[9:0] T2498;
  wire[6:0] T6072;
  wire T6073;
  wire T2499;
  wire T2500;
  wire[16:0] T2501;
  wire[16:0] T6074;
  wire[8:0] T2502;
  wire[8:0] T2503;
  wire[8:0] T6075;
  wire T2504;
  wire T2505;
  wire[7:0] T6076;
  wire T6077;
  wire[16:0] T2506;
  wire[16:0] T6078;
  wire[8:0] T2507;
  wire[7:0] T6079;
  wire T6080;
  wire T2508;
  wire T2509;
  wire[16:0] T2510;
  wire[16:0] T6081;
  wire[7:0] T2511;
  wire[7:0] T2512;
  wire[7:0] T6082;
  wire T2513;
  wire T2514;
  wire[8:0] T6083;
  wire T6084;
  wire[16:0] T2515;
  wire[16:0] T6085;
  wire[7:0] T2516;
  wire[8:0] T6086;
  wire T6087;
  wire T2517;
  wire T2518;
  wire[16:0] T2519;
  wire[16:0] T6088;
  wire[6:0] T2520;
  wire[6:0] T2521;
  wire[6:0] T6089;
  wire T2522;
  wire T2523;
  wire[9:0] T6090;
  wire T6091;
  wire[16:0] T2524;
  wire[16:0] T6092;
  wire[6:0] T2525;
  wire[9:0] T6093;
  wire T6094;
  wire T2526;
  wire T2527;
  wire[16:0] T2528;
  wire[16:0] T6095;
  wire[5:0] T2529;
  wire[5:0] T2530;
  wire[5:0] T6096;
  wire T2531;
  wire T2532;
  wire[10:0] T6097;
  wire T6098;
  wire[16:0] T2533;
  wire[16:0] T6099;
  wire[5:0] T2534;
  wire[10:0] T6100;
  wire T6101;
  wire T2535;
  wire T2536;
  wire[16:0] T2537;
  wire[16:0] T6102;
  wire[4:0] T2538;
  wire[4:0] T2539;
  wire[4:0] T6103;
  wire T2540;
  wire T2541;
  wire[11:0] T6104;
  wire T6105;
  wire[16:0] T2542;
  wire[16:0] T6106;
  wire[4:0] T2543;
  wire[11:0] T6107;
  wire T6108;
  wire T2544;
  wire T2545;
  wire[16:0] T2546;
  wire[16:0] T6109;
  wire[3:0] T2547;
  wire[3:0] T2548;
  wire[3:0] T6110;
  wire T2549;
  wire T2550;
  wire[12:0] T6111;
  wire T6112;
  wire[16:0] T2551;
  wire[16:0] T6113;
  wire[3:0] T2552;
  wire[12:0] T6114;
  wire T6115;
  wire T2553;
  wire T2554;
  wire[16:0] T2555;
  wire[16:0] T6116;
  wire[2:0] T2556;
  wire[2:0] T2557;
  wire[2:0] T6117;
  wire T2558;
  wire T2559;
  wire[13:0] T6118;
  wire T6119;
  wire[16:0] T2560;
  wire[16:0] T6120;
  wire[2:0] T2561;
  wire[13:0] T6121;
  wire T6122;
  wire T2562;
  wire T2563;
  wire[16:0] T2564;
  wire[16:0] T6123;
  wire[1:0] T2565;
  wire[1:0] T2566;
  wire[1:0] T6124;
  wire T2567;
  wire T2568;
  wire[14:0] T6125;
  wire T6126;
  wire[16:0] T2569;
  wire[16:0] T6127;
  wire[1:0] T2570;
  wire[14:0] T6128;
  wire T6129;
  wire T2571;
  wire T2572;
  wire[15:0] V_wire_en_8;
  wire[15:0] T6130;
  wire[16:0] T2573;
  wire[16:0] T2574;
  wire[16:0] T2575;
  wire[16:0] T2576;
  wire[16:0] T2577;
  wire[16:0] T2578;
  wire[16:0] T2579;
  wire[16:0] T2580;
  wire[16:0] T2581;
  wire[16:0] T2582;
  wire[16:0] T2583;
  wire[16:0] T2584;
  wire[16:0] T2585;
  wire[16:0] T2586;
  wire[16:0] T2587;
  wire[16:0] T2588;
  wire[16:0] T2589;
  wire[16:0] T2590;
  wire[16:0] T2591;
  wire[16:0] T6131;
  wire T2592;
  wire T2593;
  wire[16:0] T2594;
  wire[16:0] T2595;
  wire T2596;
  wire T2597;
  wire[3:0] T2598;
  wire T2599;
  wire T2600;
  wire[16:0] T2601;
  wire[16:0] T6132;
  wire[15:0] T2602;
  wire[15:0] T2603;
  wire[15:0] T6133;
  wire T2604;
  wire T2605;
  wire T6134;
  wire[16:0] T2606;
  wire[16:0] T6135;
  wire[15:0] T2607;
  wire T6136;
  wire T2608;
  wire T2609;
  wire[16:0] T2610;
  wire[16:0] T6137;
  wire[14:0] T2611;
  wire[14:0] T2612;
  wire[14:0] T6138;
  wire T2613;
  wire T2614;
  wire[1:0] T6139;
  wire T6140;
  wire[16:0] T2615;
  wire[16:0] T6141;
  wire[14:0] T2616;
  wire[1:0] T6142;
  wire T6143;
  wire T2617;
  wire T2618;
  wire[16:0] T2619;
  wire[16:0] T6144;
  wire[13:0] T2620;
  wire[13:0] T2621;
  wire[13:0] T6145;
  wire T2622;
  wire T2623;
  wire[2:0] T6146;
  wire T6147;
  wire[16:0] T2624;
  wire[16:0] T6148;
  wire[13:0] T2625;
  wire[2:0] T6149;
  wire T6150;
  wire T2626;
  wire T2627;
  wire[16:0] T2628;
  wire[16:0] T6151;
  wire[12:0] T2629;
  wire[12:0] T2630;
  wire[12:0] T6152;
  wire T2631;
  wire T2632;
  wire[3:0] T6153;
  wire T6154;
  wire[16:0] T2633;
  wire[16:0] T6155;
  wire[12:0] T2634;
  wire[3:0] T6156;
  wire T6157;
  wire T2635;
  wire T2636;
  wire[16:0] T2637;
  wire[16:0] T6158;
  wire[11:0] T2638;
  wire[11:0] T2639;
  wire[11:0] T6159;
  wire T2640;
  wire T2641;
  wire[4:0] T6160;
  wire T6161;
  wire[16:0] T2642;
  wire[16:0] T6162;
  wire[11:0] T2643;
  wire[4:0] T6163;
  wire T6164;
  wire T2644;
  wire T2645;
  wire[16:0] T2646;
  wire[16:0] T6165;
  wire[10:0] T2647;
  wire[10:0] T2648;
  wire[10:0] T6166;
  wire T2649;
  wire T2650;
  wire[5:0] T6167;
  wire T6168;
  wire[16:0] T2651;
  wire[16:0] T6169;
  wire[10:0] T2652;
  wire[5:0] T6170;
  wire T6171;
  wire T2653;
  wire T2654;
  wire[16:0] T2655;
  wire[16:0] T6172;
  wire[9:0] T2656;
  wire[9:0] T2657;
  wire[9:0] T6173;
  wire T2658;
  wire T2659;
  wire[6:0] T6174;
  wire T6175;
  wire[16:0] T2660;
  wire[16:0] T6176;
  wire[9:0] T2661;
  wire[6:0] T6177;
  wire T6178;
  wire T2662;
  wire T2663;
  wire[16:0] T2664;
  wire[16:0] T6179;
  wire[8:0] T2665;
  wire[8:0] T2666;
  wire[8:0] T6180;
  wire T2667;
  wire T2668;
  wire[7:0] T6181;
  wire T6182;
  wire[16:0] T2669;
  wire[16:0] T6183;
  wire[8:0] T2670;
  wire[7:0] T6184;
  wire T6185;
  wire T2671;
  wire T2672;
  wire[16:0] T2673;
  wire[16:0] T6186;
  wire[7:0] T2674;
  wire[7:0] T2675;
  wire[7:0] T6187;
  wire T2676;
  wire T2677;
  wire[8:0] T6188;
  wire T6189;
  wire[16:0] T2678;
  wire[16:0] T6190;
  wire[7:0] T2679;
  wire[8:0] T6191;
  wire T6192;
  wire T2680;
  wire T2681;
  wire[16:0] T2682;
  wire[16:0] T6193;
  wire[6:0] T2683;
  wire[6:0] T2684;
  wire[6:0] T6194;
  wire T2685;
  wire T2686;
  wire[9:0] T6195;
  wire T6196;
  wire[16:0] T2687;
  wire[16:0] T6197;
  wire[6:0] T2688;
  wire[9:0] T6198;
  wire T6199;
  wire T2689;
  wire T2690;
  wire[16:0] T2691;
  wire[16:0] T6200;
  wire[5:0] T2692;
  wire[5:0] T2693;
  wire[5:0] T6201;
  wire T2694;
  wire T2695;
  wire[10:0] T6202;
  wire T6203;
  wire[16:0] T2696;
  wire[16:0] T6204;
  wire[5:0] T2697;
  wire[10:0] T6205;
  wire T6206;
  wire T2698;
  wire T2699;
  wire[16:0] T2700;
  wire[16:0] T6207;
  wire[4:0] T2701;
  wire[4:0] T2702;
  wire[4:0] T6208;
  wire T2703;
  wire T2704;
  wire[11:0] T6209;
  wire T6210;
  wire[16:0] T2705;
  wire[16:0] T6211;
  wire[4:0] T2706;
  wire[11:0] T6212;
  wire T6213;
  wire T2707;
  wire T2708;
  wire[16:0] T2709;
  wire[16:0] T6214;
  wire[3:0] T2710;
  wire[3:0] T2711;
  wire[3:0] T6215;
  wire T2712;
  wire T2713;
  wire[12:0] T6216;
  wire T6217;
  wire[16:0] T2714;
  wire[16:0] T6218;
  wire[3:0] T2715;
  wire[12:0] T6219;
  wire T6220;
  wire T2716;
  wire T2717;
  wire[16:0] T2718;
  wire[16:0] T6221;
  wire[2:0] T2719;
  wire[2:0] T2720;
  wire[2:0] T6222;
  wire T2721;
  wire T2722;
  wire[13:0] T6223;
  wire T6224;
  wire[16:0] T2723;
  wire[16:0] T6225;
  wire[2:0] T2724;
  wire[13:0] T6226;
  wire T6227;
  wire T2725;
  wire T2726;
  wire[16:0] T2727;
  wire[16:0] T6228;
  wire[1:0] T2728;
  wire[1:0] T2729;
  wire[1:0] T6229;
  wire T2730;
  wire T2731;
  wire[14:0] T6230;
  wire T6231;
  wire[16:0] T2732;
  wire[16:0] T6232;
  wire[1:0] T2733;
  wire[14:0] T6233;
  wire T6234;
  wire T2734;
  wire T2735;
  wire[15:0] V_wire_en_9;
  wire[15:0] T6235;
  wire[16:0] T2736;
  wire[16:0] T2737;
  wire[16:0] T2738;
  wire[16:0] T2739;
  wire[16:0] T2740;
  wire[16:0] T2741;
  wire[16:0] T2742;
  wire[16:0] T2743;
  wire[16:0] T2744;
  wire[16:0] T2745;
  wire[16:0] T2746;
  wire[16:0] T2747;
  wire[16:0] T2748;
  wire[16:0] T2749;
  wire[16:0] T2750;
  wire[16:0] T2751;
  wire[16:0] T2752;
  wire[16:0] T2753;
  wire[16:0] T2754;
  wire[16:0] T6236;
  wire T2755;
  wire T2756;
  wire[16:0] T2757;
  wire[16:0] T2758;
  wire T2759;
  wire T2760;
  wire[3:0] T2761;
  wire T2762;
  wire T2763;
  wire[16:0] T2764;
  wire[16:0] T6237;
  wire[15:0] T2765;
  wire[15:0] T2766;
  wire[15:0] T6238;
  wire T2767;
  wire T2768;
  wire T6239;
  wire[16:0] T2769;
  wire[16:0] T6240;
  wire[15:0] T2770;
  wire T6241;
  wire T2771;
  wire T2772;
  wire[16:0] T2773;
  wire[16:0] T6242;
  wire[14:0] T2774;
  wire[14:0] T2775;
  wire[14:0] T6243;
  wire T2776;
  wire T2777;
  wire[1:0] T6244;
  wire T6245;
  wire[16:0] T2778;
  wire[16:0] T6246;
  wire[14:0] T2779;
  wire[1:0] T6247;
  wire T6248;
  wire T2780;
  wire T2781;
  wire[16:0] T2782;
  wire[16:0] T6249;
  wire[13:0] T2783;
  wire[13:0] T2784;
  wire[13:0] T6250;
  wire T2785;
  wire T2786;
  wire[2:0] T6251;
  wire T6252;
  wire[16:0] T2787;
  wire[16:0] T6253;
  wire[13:0] T2788;
  wire[2:0] T6254;
  wire T6255;
  wire T2789;
  wire T2790;
  wire[16:0] T2791;
  wire[16:0] T6256;
  wire[12:0] T2792;
  wire[12:0] T2793;
  wire[12:0] T6257;
  wire T2794;
  wire T2795;
  wire[3:0] T6258;
  wire T6259;
  wire[16:0] T2796;
  wire[16:0] T6260;
  wire[12:0] T2797;
  wire[3:0] T6261;
  wire T6262;
  wire T2798;
  wire T2799;
  wire[16:0] T2800;
  wire[16:0] T6263;
  wire[11:0] T2801;
  wire[11:0] T2802;
  wire[11:0] T6264;
  wire T2803;
  wire T2804;
  wire[4:0] T6265;
  wire T6266;
  wire[16:0] T2805;
  wire[16:0] T6267;
  wire[11:0] T2806;
  wire[4:0] T6268;
  wire T6269;
  wire T2807;
  wire T2808;
  wire[16:0] T2809;
  wire[16:0] T6270;
  wire[10:0] T2810;
  wire[10:0] T2811;
  wire[10:0] T6271;
  wire T2812;
  wire T2813;
  wire[5:0] T6272;
  wire T6273;
  wire[16:0] T2814;
  wire[16:0] T6274;
  wire[10:0] T2815;
  wire[5:0] T6275;
  wire T6276;
  wire T2816;
  wire T2817;
  wire[16:0] T2818;
  wire[16:0] T6277;
  wire[9:0] T2819;
  wire[9:0] T2820;
  wire[9:0] T6278;
  wire T2821;
  wire T2822;
  wire[6:0] T6279;
  wire T6280;
  wire[16:0] T2823;
  wire[16:0] T6281;
  wire[9:0] T2824;
  wire[6:0] T6282;
  wire T6283;
  wire T2825;
  wire T2826;
  wire[16:0] T2827;
  wire[16:0] T6284;
  wire[8:0] T2828;
  wire[8:0] T2829;
  wire[8:0] T6285;
  wire T2830;
  wire T2831;
  wire[7:0] T6286;
  wire T6287;
  wire[16:0] T2832;
  wire[16:0] T6288;
  wire[8:0] T2833;
  wire[7:0] T6289;
  wire T6290;
  wire T2834;
  wire T2835;
  wire[16:0] T2836;
  wire[16:0] T6291;
  wire[7:0] T2837;
  wire[7:0] T2838;
  wire[7:0] T6292;
  wire T2839;
  wire T2840;
  wire[8:0] T6293;
  wire T6294;
  wire[16:0] T2841;
  wire[16:0] T6295;
  wire[7:0] T2842;
  wire[8:0] T6296;
  wire T6297;
  wire T2843;
  wire T2844;
  wire[16:0] T2845;
  wire[16:0] T6298;
  wire[6:0] T2846;
  wire[6:0] T2847;
  wire[6:0] T6299;
  wire T2848;
  wire T2849;
  wire[9:0] T6300;
  wire T6301;
  wire[16:0] T2850;
  wire[16:0] T6302;
  wire[6:0] T2851;
  wire[9:0] T6303;
  wire T6304;
  wire T2852;
  wire T2853;
  wire[16:0] T2854;
  wire[16:0] T6305;
  wire[5:0] T2855;
  wire[5:0] T2856;
  wire[5:0] T6306;
  wire T2857;
  wire T2858;
  wire[10:0] T6307;
  wire T6308;
  wire[16:0] T2859;
  wire[16:0] T6309;
  wire[5:0] T2860;
  wire[10:0] T6310;
  wire T6311;
  wire T2861;
  wire T2862;
  wire[16:0] T2863;
  wire[16:0] T6312;
  wire[4:0] T2864;
  wire[4:0] T2865;
  wire[4:0] T6313;
  wire T2866;
  wire T2867;
  wire[11:0] T6314;
  wire T6315;
  wire[16:0] T2868;
  wire[16:0] T6316;
  wire[4:0] T2869;
  wire[11:0] T6317;
  wire T6318;
  wire T2870;
  wire T2871;
  wire[16:0] T2872;
  wire[16:0] T6319;
  wire[3:0] T2873;
  wire[3:0] T2874;
  wire[3:0] T6320;
  wire T2875;
  wire T2876;
  wire[12:0] T6321;
  wire T6322;
  wire[16:0] T2877;
  wire[16:0] T6323;
  wire[3:0] T2878;
  wire[12:0] T6324;
  wire T6325;
  wire T2879;
  wire T2880;
  wire[16:0] T2881;
  wire[16:0] T6326;
  wire[2:0] T2882;
  wire[2:0] T2883;
  wire[2:0] T6327;
  wire T2884;
  wire T2885;
  wire[13:0] T6328;
  wire T6329;
  wire[16:0] T2886;
  wire[16:0] T6330;
  wire[2:0] T2887;
  wire[13:0] T6331;
  wire T6332;
  wire T2888;
  wire T2889;
  wire[16:0] T2890;
  wire[16:0] T6333;
  wire[1:0] T2891;
  wire[1:0] T2892;
  wire[1:0] T6334;
  wire T2893;
  wire T2894;
  wire[14:0] T6335;
  wire T6336;
  wire[16:0] T2895;
  wire[16:0] T6337;
  wire[1:0] T2896;
  wire[14:0] T6338;
  wire T6339;
  wire T2897;
  wire T2898;
  wire[15:0] V_wire_en_10;
  wire[15:0] T6340;
  wire[16:0] T2899;
  wire[16:0] T2900;
  wire[16:0] T2901;
  wire[16:0] T2902;
  wire[16:0] T2903;
  wire[16:0] T2904;
  wire[16:0] T2905;
  wire[16:0] T2906;
  wire[16:0] T2907;
  wire[16:0] T2908;
  wire[16:0] T2909;
  wire[16:0] T2910;
  wire[16:0] T2911;
  wire[16:0] T2912;
  wire[16:0] T2913;
  wire[16:0] T2914;
  wire[16:0] T2915;
  wire[16:0] T2916;
  wire[16:0] T2917;
  wire[16:0] T6341;
  wire T2918;
  wire T2919;
  wire[16:0] T2920;
  wire[16:0] T2921;
  wire T2922;
  wire T2923;
  wire[3:0] T2924;
  wire T2925;
  wire T2926;
  wire[16:0] T2927;
  wire[16:0] T6342;
  wire[15:0] T2928;
  wire[15:0] T2929;
  wire[15:0] T6343;
  wire T2930;
  wire T2931;
  wire T6344;
  wire[16:0] T2932;
  wire[16:0] T6345;
  wire[15:0] T2933;
  wire T6346;
  wire T2934;
  wire T2935;
  wire[16:0] T2936;
  wire[16:0] T6347;
  wire[14:0] T2937;
  wire[14:0] T2938;
  wire[14:0] T6348;
  wire T2939;
  wire T2940;
  wire[1:0] T6349;
  wire T6350;
  wire[16:0] T2941;
  wire[16:0] T6351;
  wire[14:0] T2942;
  wire[1:0] T6352;
  wire T6353;
  wire T2943;
  wire T2944;
  wire[16:0] T2945;
  wire[16:0] T6354;
  wire[13:0] T2946;
  wire[13:0] T2947;
  wire[13:0] T6355;
  wire T2948;
  wire T2949;
  wire[2:0] T6356;
  wire T6357;
  wire[16:0] T2950;
  wire[16:0] T6358;
  wire[13:0] T2951;
  wire[2:0] T6359;
  wire T6360;
  wire T2952;
  wire T2953;
  wire[16:0] T2954;
  wire[16:0] T6361;
  wire[12:0] T2955;
  wire[12:0] T2956;
  wire[12:0] T6362;
  wire T2957;
  wire T2958;
  wire[3:0] T6363;
  wire T6364;
  wire[16:0] T2959;
  wire[16:0] T6365;
  wire[12:0] T2960;
  wire[3:0] T6366;
  wire T6367;
  wire T2961;
  wire T2962;
  wire[16:0] T2963;
  wire[16:0] T6368;
  wire[11:0] T2964;
  wire[11:0] T2965;
  wire[11:0] T6369;
  wire T2966;
  wire T2967;
  wire[4:0] T6370;
  wire T6371;
  wire[16:0] T2968;
  wire[16:0] T6372;
  wire[11:0] T2969;
  wire[4:0] T6373;
  wire T6374;
  wire T2970;
  wire T2971;
  wire[16:0] T2972;
  wire[16:0] T6375;
  wire[10:0] T2973;
  wire[10:0] T2974;
  wire[10:0] T6376;
  wire T2975;
  wire T2976;
  wire[5:0] T6377;
  wire T6378;
  wire[16:0] T2977;
  wire[16:0] T6379;
  wire[10:0] T2978;
  wire[5:0] T6380;
  wire T6381;
  wire T2979;
  wire T2980;
  wire[16:0] T2981;
  wire[16:0] T6382;
  wire[9:0] T2982;
  wire[9:0] T2983;
  wire[9:0] T6383;
  wire T2984;
  wire T2985;
  wire[6:0] T6384;
  wire T6385;
  wire[16:0] T2986;
  wire[16:0] T6386;
  wire[9:0] T2987;
  wire[6:0] T6387;
  wire T6388;
  wire T2988;
  wire T2989;
  wire[16:0] T2990;
  wire[16:0] T6389;
  wire[8:0] T2991;
  wire[8:0] T2992;
  wire[8:0] T6390;
  wire T2993;
  wire T2994;
  wire[7:0] T6391;
  wire T6392;
  wire[16:0] T2995;
  wire[16:0] T6393;
  wire[8:0] T2996;
  wire[7:0] T6394;
  wire T6395;
  wire T2997;
  wire T2998;
  wire[16:0] T2999;
  wire[16:0] T6396;
  wire[7:0] T3000;
  wire[7:0] T3001;
  wire[7:0] T6397;
  wire T3002;
  wire T3003;
  wire[8:0] T6398;
  wire T6399;
  wire[16:0] T3004;
  wire[16:0] T6400;
  wire[7:0] T3005;
  wire[8:0] T6401;
  wire T6402;
  wire T3006;
  wire T3007;
  wire[16:0] T3008;
  wire[16:0] T6403;
  wire[6:0] T3009;
  wire[6:0] T3010;
  wire[6:0] T6404;
  wire T3011;
  wire T3012;
  wire[9:0] T6405;
  wire T6406;
  wire[16:0] T3013;
  wire[16:0] T6407;
  wire[6:0] T3014;
  wire[9:0] T6408;
  wire T6409;
  wire T3015;
  wire T3016;
  wire[16:0] T3017;
  wire[16:0] T6410;
  wire[5:0] T3018;
  wire[5:0] T3019;
  wire[5:0] T6411;
  wire T3020;
  wire T3021;
  wire[10:0] T6412;
  wire T6413;
  wire[16:0] T3022;
  wire[16:0] T6414;
  wire[5:0] T3023;
  wire[10:0] T6415;
  wire T6416;
  wire T3024;
  wire T3025;
  wire[16:0] T3026;
  wire[16:0] T6417;
  wire[4:0] T3027;
  wire[4:0] T3028;
  wire[4:0] T6418;
  wire T3029;
  wire T3030;
  wire[11:0] T6419;
  wire T6420;
  wire[16:0] T3031;
  wire[16:0] T6421;
  wire[4:0] T3032;
  wire[11:0] T6422;
  wire T6423;
  wire T3033;
  wire T3034;
  wire[16:0] T3035;
  wire[16:0] T6424;
  wire[3:0] T3036;
  wire[3:0] T3037;
  wire[3:0] T6425;
  wire T3038;
  wire T3039;
  wire[12:0] T6426;
  wire T6427;
  wire[16:0] T3040;
  wire[16:0] T6428;
  wire[3:0] T3041;
  wire[12:0] T6429;
  wire T6430;
  wire T3042;
  wire T3043;
  wire[16:0] T3044;
  wire[16:0] T6431;
  wire[2:0] T3045;
  wire[2:0] T3046;
  wire[2:0] T6432;
  wire T3047;
  wire T3048;
  wire[13:0] T6433;
  wire T6434;
  wire[16:0] T3049;
  wire[16:0] T6435;
  wire[2:0] T3050;
  wire[13:0] T6436;
  wire T6437;
  wire T3051;
  wire T3052;
  wire[16:0] T3053;
  wire[16:0] T6438;
  wire[1:0] T3054;
  wire[1:0] T3055;
  wire[1:0] T6439;
  wire T3056;
  wire T3057;
  wire[14:0] T6440;
  wire T6441;
  wire[16:0] T3058;
  wire[16:0] T6442;
  wire[1:0] T3059;
  wire[14:0] T6443;
  wire T6444;
  wire T3060;
  wire T3061;
  wire[15:0] V_wire_en_11;
  wire[15:0] T6445;
  wire[16:0] T3062;
  wire[16:0] T3063;
  wire[16:0] T3064;
  wire[16:0] T3065;
  wire[16:0] T3066;
  wire[16:0] T3067;
  wire[16:0] T3068;
  wire[16:0] T3069;
  wire[16:0] T3070;
  wire[16:0] T3071;
  wire[16:0] T3072;
  wire[16:0] T3073;
  wire[16:0] T3074;
  wire[16:0] T3075;
  wire[16:0] T3076;
  wire[16:0] T3077;
  wire[16:0] T3078;
  wire[16:0] T3079;
  wire[16:0] T3080;
  wire[16:0] T6446;
  wire T3081;
  wire T3082;
  wire[16:0] T3083;
  wire[16:0] T3084;
  wire T3085;
  wire T3086;
  wire[3:0] T3087;
  wire T3088;
  wire T3089;
  wire[16:0] T3090;
  wire[16:0] T6447;
  wire[15:0] T3091;
  wire[15:0] T3092;
  wire[15:0] T6448;
  wire T3093;
  wire T3094;
  wire T6449;
  wire[16:0] T3095;
  wire[16:0] T6450;
  wire[15:0] T3096;
  wire T6451;
  wire T3097;
  wire T3098;
  wire[16:0] T3099;
  wire[16:0] T6452;
  wire[14:0] T3100;
  wire[14:0] T3101;
  wire[14:0] T6453;
  wire T3102;
  wire T3103;
  wire[1:0] T6454;
  wire T6455;
  wire[16:0] T3104;
  wire[16:0] T6456;
  wire[14:0] T3105;
  wire[1:0] T6457;
  wire T6458;
  wire T3106;
  wire T3107;
  wire[16:0] T3108;
  wire[16:0] T6459;
  wire[13:0] T3109;
  wire[13:0] T3110;
  wire[13:0] T6460;
  wire T3111;
  wire T3112;
  wire[2:0] T6461;
  wire T6462;
  wire[16:0] T3113;
  wire[16:0] T6463;
  wire[13:0] T3114;
  wire[2:0] T6464;
  wire T6465;
  wire T3115;
  wire T3116;
  wire[16:0] T3117;
  wire[16:0] T6466;
  wire[12:0] T3118;
  wire[12:0] T3119;
  wire[12:0] T6467;
  wire T3120;
  wire T3121;
  wire[3:0] T6468;
  wire T6469;
  wire[16:0] T3122;
  wire[16:0] T6470;
  wire[12:0] T3123;
  wire[3:0] T6471;
  wire T6472;
  wire T3124;
  wire T3125;
  wire[16:0] T3126;
  wire[16:0] T6473;
  wire[11:0] T3127;
  wire[11:0] T3128;
  wire[11:0] T6474;
  wire T3129;
  wire T3130;
  wire[4:0] T6475;
  wire T6476;
  wire[16:0] T3131;
  wire[16:0] T6477;
  wire[11:0] T3132;
  wire[4:0] T6478;
  wire T6479;
  wire T3133;
  wire T3134;
  wire[16:0] T3135;
  wire[16:0] T6480;
  wire[10:0] T3136;
  wire[10:0] T3137;
  wire[10:0] T6481;
  wire T3138;
  wire T3139;
  wire[5:0] T6482;
  wire T6483;
  wire[16:0] T3140;
  wire[16:0] T6484;
  wire[10:0] T3141;
  wire[5:0] T6485;
  wire T6486;
  wire T3142;
  wire T3143;
  wire[16:0] T3144;
  wire[16:0] T6487;
  wire[9:0] T3145;
  wire[9:0] T3146;
  wire[9:0] T6488;
  wire T3147;
  wire T3148;
  wire[6:0] T6489;
  wire T6490;
  wire[16:0] T3149;
  wire[16:0] T6491;
  wire[9:0] T3150;
  wire[6:0] T6492;
  wire T6493;
  wire T3151;
  wire T3152;
  wire[16:0] T3153;
  wire[16:0] T6494;
  wire[8:0] T3154;
  wire[8:0] T3155;
  wire[8:0] T6495;
  wire T3156;
  wire T3157;
  wire[7:0] T6496;
  wire T6497;
  wire[16:0] T3158;
  wire[16:0] T6498;
  wire[8:0] T3159;
  wire[7:0] T6499;
  wire T6500;
  wire T3160;
  wire T3161;
  wire[16:0] T3162;
  wire[16:0] T6501;
  wire[7:0] T3163;
  wire[7:0] T3164;
  wire[7:0] T6502;
  wire T3165;
  wire T3166;
  wire[8:0] T6503;
  wire T6504;
  wire[16:0] T3167;
  wire[16:0] T6505;
  wire[7:0] T3168;
  wire[8:0] T6506;
  wire T6507;
  wire T3169;
  wire T3170;
  wire[16:0] T3171;
  wire[16:0] T6508;
  wire[6:0] T3172;
  wire[6:0] T3173;
  wire[6:0] T6509;
  wire T3174;
  wire T3175;
  wire[9:0] T6510;
  wire T6511;
  wire[16:0] T3176;
  wire[16:0] T6512;
  wire[6:0] T3177;
  wire[9:0] T6513;
  wire T6514;
  wire T3178;
  wire T3179;
  wire[16:0] T3180;
  wire[16:0] T6515;
  wire[5:0] T3181;
  wire[5:0] T3182;
  wire[5:0] T6516;
  wire T3183;
  wire T3184;
  wire[10:0] T6517;
  wire T6518;
  wire[16:0] T3185;
  wire[16:0] T6519;
  wire[5:0] T3186;
  wire[10:0] T6520;
  wire T6521;
  wire T3187;
  wire T3188;
  wire[16:0] T3189;
  wire[16:0] T6522;
  wire[4:0] T3190;
  wire[4:0] T3191;
  wire[4:0] T6523;
  wire T3192;
  wire T3193;
  wire[11:0] T6524;
  wire T6525;
  wire[16:0] T3194;
  wire[16:0] T6526;
  wire[4:0] T3195;
  wire[11:0] T6527;
  wire T6528;
  wire T3196;
  wire T3197;
  wire[16:0] T3198;
  wire[16:0] T6529;
  wire[3:0] T3199;
  wire[3:0] T3200;
  wire[3:0] T6530;
  wire T3201;
  wire T3202;
  wire[12:0] T6531;
  wire T6532;
  wire[16:0] T3203;
  wire[16:0] T6533;
  wire[3:0] T3204;
  wire[12:0] T6534;
  wire T6535;
  wire T3205;
  wire T3206;
  wire[16:0] T3207;
  wire[16:0] T6536;
  wire[2:0] T3208;
  wire[2:0] T3209;
  wire[2:0] T6537;
  wire T3210;
  wire T3211;
  wire[13:0] T6538;
  wire T6539;
  wire[16:0] T3212;
  wire[16:0] T6540;
  wire[2:0] T3213;
  wire[13:0] T6541;
  wire T6542;
  wire T3214;
  wire T3215;
  wire[16:0] T3216;
  wire[16:0] T6543;
  wire[1:0] T3217;
  wire[1:0] T3218;
  wire[1:0] T6544;
  wire T3219;
  wire T3220;
  wire[14:0] T6545;
  wire T6546;
  wire[16:0] T3221;
  wire[16:0] T6547;
  wire[1:0] T3222;
  wire[14:0] T6548;
  wire T6549;
  wire T3223;
  wire T3224;
  wire[15:0] V_wire_en_12;
  wire[15:0] T6550;
  wire[16:0] T3225;
  wire[16:0] T3226;
  wire[16:0] T3227;
  wire[16:0] T3228;
  wire[16:0] T3229;
  wire[16:0] T3230;
  wire[16:0] T3231;
  wire[16:0] T3232;
  wire[16:0] T3233;
  wire[16:0] T3234;
  wire[16:0] T3235;
  wire[16:0] T3236;
  wire[16:0] T3237;
  wire[16:0] T3238;
  wire[16:0] T3239;
  wire[16:0] T3240;
  wire[16:0] T3241;
  wire[16:0] T3242;
  wire[16:0] T3243;
  wire[16:0] T6551;
  wire T3244;
  wire T3245;
  wire[16:0] T3246;
  wire[16:0] T3247;
  wire T3248;
  wire T3249;
  wire[3:0] T3250;
  wire T3251;
  wire T3252;
  wire[16:0] T3253;
  wire[16:0] T6552;
  wire[15:0] T3254;
  wire[15:0] T3255;
  wire[15:0] T6553;
  wire T3256;
  wire T3257;
  wire T6554;
  wire[16:0] T3258;
  wire[16:0] T6555;
  wire[15:0] T3259;
  wire T6556;
  wire T3260;
  wire T3261;
  wire[16:0] T3262;
  wire[16:0] T6557;
  wire[14:0] T3263;
  wire[14:0] T3264;
  wire[14:0] T6558;
  wire T3265;
  wire T3266;
  wire[1:0] T6559;
  wire T6560;
  wire[16:0] T3267;
  wire[16:0] T6561;
  wire[14:0] T3268;
  wire[1:0] T6562;
  wire T6563;
  wire T3269;
  wire T3270;
  wire[16:0] T3271;
  wire[16:0] T6564;
  wire[13:0] T3272;
  wire[13:0] T3273;
  wire[13:0] T6565;
  wire T3274;
  wire T3275;
  wire[2:0] T6566;
  wire T6567;
  wire[16:0] T3276;
  wire[16:0] T6568;
  wire[13:0] T3277;
  wire[2:0] T6569;
  wire T6570;
  wire T3278;
  wire T3279;
  wire[16:0] T3280;
  wire[16:0] T6571;
  wire[12:0] T3281;
  wire[12:0] T3282;
  wire[12:0] T6572;
  wire T3283;
  wire T3284;
  wire[3:0] T6573;
  wire T6574;
  wire[16:0] T3285;
  wire[16:0] T6575;
  wire[12:0] T3286;
  wire[3:0] T6576;
  wire T6577;
  wire T3287;
  wire T3288;
  wire[16:0] T3289;
  wire[16:0] T6578;
  wire[11:0] T3290;
  wire[11:0] T3291;
  wire[11:0] T6579;
  wire T3292;
  wire T3293;
  wire[4:0] T6580;
  wire T6581;
  wire[16:0] T3294;
  wire[16:0] T6582;
  wire[11:0] T3295;
  wire[4:0] T6583;
  wire T6584;
  wire T3296;
  wire T3297;
  wire[16:0] T3298;
  wire[16:0] T6585;
  wire[10:0] T3299;
  wire[10:0] T3300;
  wire[10:0] T6586;
  wire T3301;
  wire T3302;
  wire[5:0] T6587;
  wire T6588;
  wire[16:0] T3303;
  wire[16:0] T6589;
  wire[10:0] T3304;
  wire[5:0] T6590;
  wire T6591;
  wire T3305;
  wire T3306;
  wire[16:0] T3307;
  wire[16:0] T6592;
  wire[9:0] T3308;
  wire[9:0] T3309;
  wire[9:0] T6593;
  wire T3310;
  wire T3311;
  wire[6:0] T6594;
  wire T6595;
  wire[16:0] T3312;
  wire[16:0] T6596;
  wire[9:0] T3313;
  wire[6:0] T6597;
  wire T6598;
  wire T3314;
  wire T3315;
  wire[16:0] T3316;
  wire[16:0] T6599;
  wire[8:0] T3317;
  wire[8:0] T3318;
  wire[8:0] T6600;
  wire T3319;
  wire T3320;
  wire[7:0] T6601;
  wire T6602;
  wire[16:0] T3321;
  wire[16:0] T6603;
  wire[8:0] T3322;
  wire[7:0] T6604;
  wire T6605;
  wire T3323;
  wire T3324;
  wire[16:0] T3325;
  wire[16:0] T6606;
  wire[7:0] T3326;
  wire[7:0] T3327;
  wire[7:0] T6607;
  wire T3328;
  wire T3329;
  wire[8:0] T6608;
  wire T6609;
  wire[16:0] T3330;
  wire[16:0] T6610;
  wire[7:0] T3331;
  wire[8:0] T6611;
  wire T6612;
  wire T3332;
  wire T3333;
  wire[16:0] T3334;
  wire[16:0] T6613;
  wire[6:0] T3335;
  wire[6:0] T3336;
  wire[6:0] T6614;
  wire T3337;
  wire T3338;
  wire[9:0] T6615;
  wire T6616;
  wire[16:0] T3339;
  wire[16:0] T6617;
  wire[6:0] T3340;
  wire[9:0] T6618;
  wire T6619;
  wire T3341;
  wire T3342;
  wire[16:0] T3343;
  wire[16:0] T6620;
  wire[5:0] T3344;
  wire[5:0] T3345;
  wire[5:0] T6621;
  wire T3346;
  wire T3347;
  wire[10:0] T6622;
  wire T6623;
  wire[16:0] T3348;
  wire[16:0] T6624;
  wire[5:0] T3349;
  wire[10:0] T6625;
  wire T6626;
  wire T3350;
  wire T3351;
  wire[16:0] T3352;
  wire[16:0] T6627;
  wire[4:0] T3353;
  wire[4:0] T3354;
  wire[4:0] T6628;
  wire T3355;
  wire T3356;
  wire[11:0] T6629;
  wire T6630;
  wire[16:0] T3357;
  wire[16:0] T6631;
  wire[4:0] T3358;
  wire[11:0] T6632;
  wire T6633;
  wire T3359;
  wire T3360;
  wire[16:0] T3361;
  wire[16:0] T6634;
  wire[3:0] T3362;
  wire[3:0] T3363;
  wire[3:0] T6635;
  wire T3364;
  wire T3365;
  wire[12:0] T6636;
  wire T6637;
  wire[16:0] T3366;
  wire[16:0] T6638;
  wire[3:0] T3367;
  wire[12:0] T6639;
  wire T6640;
  wire T3368;
  wire T3369;
  wire[16:0] T3370;
  wire[16:0] T6641;
  wire[2:0] T3371;
  wire[2:0] T3372;
  wire[2:0] T6642;
  wire T3373;
  wire T3374;
  wire[13:0] T6643;
  wire T6644;
  wire[16:0] T3375;
  wire[16:0] T6645;
  wire[2:0] T3376;
  wire[13:0] T6646;
  wire T6647;
  wire T3377;
  wire T3378;
  wire[16:0] T3379;
  wire[16:0] T6648;
  wire[1:0] T3380;
  wire[1:0] T3381;
  wire[1:0] T6649;
  wire T3382;
  wire T3383;
  wire[14:0] T6650;
  wire T6651;
  wire[16:0] T3384;
  wire[16:0] T6652;
  wire[1:0] T3385;
  wire[14:0] T6653;
  wire T6654;
  wire T3386;
  wire T3387;
  wire[15:0] V_wire_en_13;
  wire[15:0] T6655;
  wire[16:0] T3388;
  wire[16:0] T3389;
  wire[16:0] T3390;
  wire[16:0] T3391;
  wire[16:0] T3392;
  wire[16:0] T3393;
  wire[16:0] T3394;
  wire[16:0] T3395;
  wire[16:0] T3396;
  wire[16:0] T3397;
  wire[16:0] T3398;
  wire[16:0] T3399;
  wire[16:0] T3400;
  wire[16:0] T3401;
  wire[16:0] T3402;
  wire[16:0] T3403;
  wire[16:0] T3404;
  wire[16:0] T3405;
  wire[16:0] T3406;
  wire[16:0] T6656;
  wire T3407;
  wire T3408;
  wire[16:0] T3409;
  wire[16:0] T3410;
  wire T3411;
  wire T3412;
  wire[3:0] T3413;
  wire T3414;
  wire T3415;
  wire[16:0] T3416;
  wire[16:0] T6657;
  wire[15:0] T3417;
  wire[15:0] T3418;
  wire[15:0] T6658;
  wire T3419;
  wire T3420;
  wire T6659;
  wire[16:0] T3421;
  wire[16:0] T6660;
  wire[15:0] T3422;
  wire T6661;
  wire T3423;
  wire T3424;
  wire[16:0] T3425;
  wire[16:0] T6662;
  wire[14:0] T3426;
  wire[14:0] T3427;
  wire[14:0] T6663;
  wire T3428;
  wire T3429;
  wire[1:0] T6664;
  wire T6665;
  wire[16:0] T3430;
  wire[16:0] T6666;
  wire[14:0] T3431;
  wire[1:0] T6667;
  wire T6668;
  wire T3432;
  wire T3433;
  wire[16:0] T3434;
  wire[16:0] T6669;
  wire[13:0] T3435;
  wire[13:0] T3436;
  wire[13:0] T6670;
  wire T3437;
  wire T3438;
  wire[2:0] T6671;
  wire T6672;
  wire[16:0] T3439;
  wire[16:0] T6673;
  wire[13:0] T3440;
  wire[2:0] T6674;
  wire T6675;
  wire T3441;
  wire T3442;
  wire[16:0] T3443;
  wire[16:0] T6676;
  wire[12:0] T3444;
  wire[12:0] T3445;
  wire[12:0] T6677;
  wire T3446;
  wire T3447;
  wire[3:0] T6678;
  wire T6679;
  wire[16:0] T3448;
  wire[16:0] T6680;
  wire[12:0] T3449;
  wire[3:0] T6681;
  wire T6682;
  wire T3450;
  wire T3451;
  wire[16:0] T3452;
  wire[16:0] T6683;
  wire[11:0] T3453;
  wire[11:0] T3454;
  wire[11:0] T6684;
  wire T3455;
  wire T3456;
  wire[4:0] T6685;
  wire T6686;
  wire[16:0] T3457;
  wire[16:0] T6687;
  wire[11:0] T3458;
  wire[4:0] T6688;
  wire T6689;
  wire T3459;
  wire T3460;
  wire[16:0] T3461;
  wire[16:0] T6690;
  wire[10:0] T3462;
  wire[10:0] T3463;
  wire[10:0] T6691;
  wire T3464;
  wire T3465;
  wire[5:0] T6692;
  wire T6693;
  wire[16:0] T3466;
  wire[16:0] T6694;
  wire[10:0] T3467;
  wire[5:0] T6695;
  wire T6696;
  wire T3468;
  wire T3469;
  wire[16:0] T3470;
  wire[16:0] T6697;
  wire[9:0] T3471;
  wire[9:0] T3472;
  wire[9:0] T6698;
  wire T3473;
  wire T3474;
  wire[6:0] T6699;
  wire T6700;
  wire[16:0] T3475;
  wire[16:0] T6701;
  wire[9:0] T3476;
  wire[6:0] T6702;
  wire T6703;
  wire T3477;
  wire T3478;
  wire[16:0] T3479;
  wire[16:0] T6704;
  wire[8:0] T3480;
  wire[8:0] T3481;
  wire[8:0] T6705;
  wire T3482;
  wire T3483;
  wire[7:0] T6706;
  wire T6707;
  wire[16:0] T3484;
  wire[16:0] T6708;
  wire[8:0] T3485;
  wire[7:0] T6709;
  wire T6710;
  wire T3486;
  wire T3487;
  wire[16:0] T3488;
  wire[16:0] T6711;
  wire[7:0] T3489;
  wire[7:0] T3490;
  wire[7:0] T6712;
  wire T3491;
  wire T3492;
  wire[8:0] T6713;
  wire T6714;
  wire[16:0] T3493;
  wire[16:0] T6715;
  wire[7:0] T3494;
  wire[8:0] T6716;
  wire T6717;
  wire T3495;
  wire T3496;
  wire[16:0] T3497;
  wire[16:0] T6718;
  wire[6:0] T3498;
  wire[6:0] T3499;
  wire[6:0] T6719;
  wire T3500;
  wire T3501;
  wire[9:0] T6720;
  wire T6721;
  wire[16:0] T3502;
  wire[16:0] T6722;
  wire[6:0] T3503;
  wire[9:0] T6723;
  wire T6724;
  wire T3504;
  wire T3505;
  wire[16:0] T3506;
  wire[16:0] T6725;
  wire[5:0] T3507;
  wire[5:0] T3508;
  wire[5:0] T6726;
  wire T3509;
  wire T3510;
  wire[10:0] T6727;
  wire T6728;
  wire[16:0] T3511;
  wire[16:0] T6729;
  wire[5:0] T3512;
  wire[10:0] T6730;
  wire T6731;
  wire T3513;
  wire T3514;
  wire[16:0] T3515;
  wire[16:0] T6732;
  wire[4:0] T3516;
  wire[4:0] T3517;
  wire[4:0] T6733;
  wire T3518;
  wire T3519;
  wire[11:0] T6734;
  wire T6735;
  wire[16:0] T3520;
  wire[16:0] T6736;
  wire[4:0] T3521;
  wire[11:0] T6737;
  wire T6738;
  wire T3522;
  wire T3523;
  wire[16:0] T3524;
  wire[16:0] T6739;
  wire[3:0] T3525;
  wire[3:0] T3526;
  wire[3:0] T6740;
  wire T3527;
  wire T3528;
  wire[12:0] T6741;
  wire T6742;
  wire[16:0] T3529;
  wire[16:0] T6743;
  wire[3:0] T3530;
  wire[12:0] T6744;
  wire T6745;
  wire T3531;
  wire T3532;
  wire[16:0] T3533;
  wire[16:0] T6746;
  wire[2:0] T3534;
  wire[2:0] T3535;
  wire[2:0] T6747;
  wire T3536;
  wire T3537;
  wire[13:0] T6748;
  wire T6749;
  wire[16:0] T3538;
  wire[16:0] T6750;
  wire[2:0] T3539;
  wire[13:0] T6751;
  wire T6752;
  wire T3540;
  wire T3541;
  wire[16:0] T3542;
  wire[16:0] T6753;
  wire[1:0] T3543;
  wire[1:0] T3544;
  wire[1:0] T6754;
  wire T3545;
  wire T3546;
  wire[14:0] T6755;
  wire T6756;
  wire[16:0] T3547;
  wire[16:0] T6757;
  wire[1:0] T3548;
  wire[14:0] T6758;
  wire T6759;
  wire T3549;
  wire T3550;
  wire[15:0] V_wire_en_14;
  wire[15:0] T6760;
  wire[16:0] T3551;
  wire[16:0] T3552;
  wire[16:0] T3553;
  wire[16:0] T3554;
  wire[16:0] T3555;
  wire[16:0] T3556;
  wire[16:0] T3557;
  wire[16:0] T3558;
  wire[16:0] T3559;
  wire[16:0] T3560;
  wire[16:0] T3561;
  wire[16:0] T3562;
  wire[16:0] T3563;
  wire[16:0] T3564;
  wire[16:0] T3565;
  wire[16:0] T3566;
  wire[16:0] T3567;
  wire[16:0] T3568;
  wire[16:0] T3569;
  wire[16:0] T6761;
  wire T3570;
  wire T3571;
  wire[16:0] T3572;
  wire[16:0] T3573;
  wire T3574;
  wire T3575;
  wire[3:0] T3576;
  wire T3577;
  wire T3578;
  wire[16:0] T3579;
  wire[16:0] T6762;
  wire[15:0] T3580;
  wire[15:0] T3581;
  wire[15:0] T6763;
  wire T3582;
  wire T3583;
  wire T6764;
  wire[16:0] T3584;
  wire[16:0] T6765;
  wire[15:0] T3585;
  wire T6766;
  wire T3586;
  wire T3587;
  wire[16:0] T3588;
  wire[16:0] T6767;
  wire[14:0] T3589;
  wire[14:0] T3590;
  wire[14:0] T6768;
  wire T3591;
  wire T3592;
  wire[1:0] T6769;
  wire T6770;
  wire[16:0] T3593;
  wire[16:0] T6771;
  wire[14:0] T3594;
  wire[1:0] T6772;
  wire T6773;
  wire T3595;
  wire T3596;
  wire[16:0] T3597;
  wire[16:0] T6774;
  wire[13:0] T3598;
  wire[13:0] T3599;
  wire[13:0] T6775;
  wire T3600;
  wire T3601;
  wire[2:0] T6776;
  wire T6777;
  wire[16:0] T3602;
  wire[16:0] T6778;
  wire[13:0] T3603;
  wire[2:0] T6779;
  wire T6780;
  wire T3604;
  wire T3605;
  wire[16:0] T3606;
  wire[16:0] T6781;
  wire[12:0] T3607;
  wire[12:0] T3608;
  wire[12:0] T6782;
  wire T3609;
  wire T3610;
  wire[3:0] T6783;
  wire T6784;
  wire[16:0] T3611;
  wire[16:0] T6785;
  wire[12:0] T3612;
  wire[3:0] T6786;
  wire T6787;
  wire T3613;
  wire T3614;
  wire[16:0] T3615;
  wire[16:0] T6788;
  wire[11:0] T3616;
  wire[11:0] T3617;
  wire[11:0] T6789;
  wire T3618;
  wire T3619;
  wire[4:0] T6790;
  wire T6791;
  wire[16:0] T3620;
  wire[16:0] T6792;
  wire[11:0] T3621;
  wire[4:0] T6793;
  wire T6794;
  wire T3622;
  wire T3623;
  wire[16:0] T3624;
  wire[16:0] T6795;
  wire[10:0] T3625;
  wire[10:0] T3626;
  wire[10:0] T6796;
  wire T3627;
  wire T3628;
  wire[5:0] T6797;
  wire T6798;
  wire[16:0] T3629;
  wire[16:0] T6799;
  wire[10:0] T3630;
  wire[5:0] T6800;
  wire T6801;
  wire T3631;
  wire T3632;
  wire[16:0] T3633;
  wire[16:0] T6802;
  wire[9:0] T3634;
  wire[9:0] T3635;
  wire[9:0] T6803;
  wire T3636;
  wire T3637;
  wire[6:0] T6804;
  wire T6805;
  wire[16:0] T3638;
  wire[16:0] T6806;
  wire[9:0] T3639;
  wire[6:0] T6807;
  wire T6808;
  wire T3640;
  wire T3641;
  wire[16:0] T3642;
  wire[16:0] T6809;
  wire[8:0] T3643;
  wire[8:0] T3644;
  wire[8:0] T6810;
  wire T3645;
  wire T3646;
  wire[7:0] T6811;
  wire T6812;
  wire[16:0] T3647;
  wire[16:0] T6813;
  wire[8:0] T3648;
  wire[7:0] T6814;
  wire T6815;
  wire T3649;
  wire T3650;
  wire[16:0] T3651;
  wire[16:0] T6816;
  wire[7:0] T3652;
  wire[7:0] T3653;
  wire[7:0] T6817;
  wire T3654;
  wire T3655;
  wire[8:0] T6818;
  wire T6819;
  wire[16:0] T3656;
  wire[16:0] T6820;
  wire[7:0] T3657;
  wire[8:0] T6821;
  wire T6822;
  wire T3658;
  wire T3659;
  wire[16:0] T3660;
  wire[16:0] T6823;
  wire[6:0] T3661;
  wire[6:0] T3662;
  wire[6:0] T6824;
  wire T3663;
  wire T3664;
  wire[9:0] T6825;
  wire T6826;
  wire[16:0] T3665;
  wire[16:0] T6827;
  wire[6:0] T3666;
  wire[9:0] T6828;
  wire T6829;
  wire T3667;
  wire T3668;
  wire[16:0] T3669;
  wire[16:0] T6830;
  wire[5:0] T3670;
  wire[5:0] T3671;
  wire[5:0] T6831;
  wire T3672;
  wire T3673;
  wire[10:0] T6832;
  wire T6833;
  wire[16:0] T3674;
  wire[16:0] T6834;
  wire[5:0] T3675;
  wire[10:0] T6835;
  wire T6836;
  wire T3676;
  wire T3677;
  wire[16:0] T3678;
  wire[16:0] T6837;
  wire[4:0] T3679;
  wire[4:0] T3680;
  wire[4:0] T6838;
  wire T3681;
  wire T3682;
  wire[11:0] T6839;
  wire T6840;
  wire[16:0] T3683;
  wire[16:0] T6841;
  wire[4:0] T3684;
  wire[11:0] T6842;
  wire T6843;
  wire T3685;
  wire T3686;
  wire[16:0] T3687;
  wire[16:0] T6844;
  wire[3:0] T3688;
  wire[3:0] T3689;
  wire[3:0] T6845;
  wire T3690;
  wire T3691;
  wire[12:0] T6846;
  wire T6847;
  wire[16:0] T3692;
  wire[16:0] T6848;
  wire[3:0] T3693;
  wire[12:0] T6849;
  wire T6850;
  wire T3694;
  wire T3695;
  wire[16:0] T3696;
  wire[16:0] T6851;
  wire[2:0] T3697;
  wire[2:0] T3698;
  wire[2:0] T6852;
  wire T3699;
  wire T3700;
  wire[13:0] T6853;
  wire T6854;
  wire[16:0] T3701;
  wire[16:0] T6855;
  wire[2:0] T3702;
  wire[13:0] T6856;
  wire T6857;
  wire T3703;
  wire T3704;
  wire[16:0] T3705;
  wire[16:0] T6858;
  wire[1:0] T3706;
  wire[1:0] T3707;
  wire[1:0] T6859;
  wire T3708;
  wire T3709;
  wire[14:0] T6860;
  wire T6861;
  wire[16:0] T3710;
  wire[16:0] T6862;
  wire[1:0] T3711;
  wire[14:0] T6863;
  wire T6864;
  wire T3712;
  wire T3713;
  wire[15:0] V_wire_en_15;
  wire[15:0] T6865;
  wire[16:0] T3714;
  wire[16:0] T3715;
  wire[16:0] T3716;
  wire[16:0] T3717;
  wire[16:0] T3718;
  wire[16:0] T3719;
  wire[16:0] T3720;
  wire[16:0] T3721;
  wire[16:0] T3722;
  wire[16:0] T3723;
  wire[16:0] T3724;
  wire[16:0] T3725;
  wire[16:0] T3726;
  wire[16:0] T3727;
  wire[16:0] T3728;
  wire[16:0] T3729;
  wire[16:0] T3730;
  wire[16:0] T3731;
  wire[16:0] T3732;
  wire[16:0] T6866;
  wire T3733;
  wire T3734;
  wire[16:0] T3735;
  wire[16:0] T3736;
  wire T3737;
  wire T3738;
  wire[3:0] T3739;
  wire T3740;
  wire T3741;
  wire[16:0] T3742;
  wire[16:0] T6867;
  wire[15:0] T3743;
  wire[15:0] T3744;
  wire[15:0] T6868;
  wire T3745;
  wire T3746;
  wire T6869;
  wire[16:0] T3747;
  wire[16:0] T6870;
  wire[15:0] T3748;
  wire T6871;
  wire T3749;
  wire T3750;
  wire[16:0] T3751;
  wire[16:0] T6872;
  wire[14:0] T3752;
  wire[14:0] T3753;
  wire[14:0] T6873;
  wire T3754;
  wire T3755;
  wire[1:0] T6874;
  wire T6875;
  wire[16:0] T3756;
  wire[16:0] T6876;
  wire[14:0] T3757;
  wire[1:0] T6877;
  wire T6878;
  wire T3758;
  wire T3759;
  wire[16:0] T3760;
  wire[16:0] T6879;
  wire[13:0] T3761;
  wire[13:0] T3762;
  wire[13:0] T6880;
  wire T3763;
  wire T3764;
  wire[2:0] T6881;
  wire T6882;
  wire[16:0] T3765;
  wire[16:0] T6883;
  wire[13:0] T3766;
  wire[2:0] T6884;
  wire T6885;
  wire T3767;
  wire T3768;
  wire[16:0] T3769;
  wire[16:0] T6886;
  wire[12:0] T3770;
  wire[12:0] T3771;
  wire[12:0] T6887;
  wire T3772;
  wire T3773;
  wire[3:0] T6888;
  wire T6889;
  wire[16:0] T3774;
  wire[16:0] T6890;
  wire[12:0] T3775;
  wire[3:0] T6891;
  wire T6892;
  wire T3776;
  wire T3777;
  wire[16:0] T3778;
  wire[16:0] T6893;
  wire[11:0] T3779;
  wire[11:0] T3780;
  wire[11:0] T6894;
  wire T3781;
  wire T3782;
  wire[4:0] T6895;
  wire T6896;
  wire[16:0] T3783;
  wire[16:0] T6897;
  wire[11:0] T3784;
  wire[4:0] T6898;
  wire T6899;
  wire T3785;
  wire T3786;
  wire[16:0] T3787;
  wire[16:0] T6900;
  wire[10:0] T3788;
  wire[10:0] T3789;
  wire[10:0] T6901;
  wire T3790;
  wire T3791;
  wire[5:0] T6902;
  wire T6903;
  wire[16:0] T3792;
  wire[16:0] T6904;
  wire[10:0] T3793;
  wire[5:0] T6905;
  wire T6906;
  wire T3794;
  wire T3795;
  wire[16:0] T3796;
  wire[16:0] T6907;
  wire[9:0] T3797;
  wire[9:0] T3798;
  wire[9:0] T6908;
  wire T3799;
  wire T3800;
  wire[6:0] T6909;
  wire T6910;
  wire[16:0] T3801;
  wire[16:0] T6911;
  wire[9:0] T3802;
  wire[6:0] T6912;
  wire T6913;
  wire T3803;
  wire T3804;
  wire[16:0] T3805;
  wire[16:0] T6914;
  wire[8:0] T3806;
  wire[8:0] T3807;
  wire[8:0] T6915;
  wire T3808;
  wire T3809;
  wire[7:0] T6916;
  wire T6917;
  wire[16:0] T3810;
  wire[16:0] T6918;
  wire[8:0] T3811;
  wire[7:0] T6919;
  wire T6920;
  wire T3812;
  wire T3813;
  wire[16:0] T3814;
  wire[16:0] T6921;
  wire[7:0] T3815;
  wire[7:0] T3816;
  wire[7:0] T6922;
  wire T3817;
  wire T3818;
  wire[8:0] T6923;
  wire T6924;
  wire[16:0] T3819;
  wire[16:0] T6925;
  wire[7:0] T3820;
  wire[8:0] T6926;
  wire T6927;
  wire T3821;
  wire T3822;
  wire[16:0] T3823;
  wire[16:0] T6928;
  wire[6:0] T3824;
  wire[6:0] T3825;
  wire[6:0] T6929;
  wire T3826;
  wire T3827;
  wire[9:0] T6930;
  wire T6931;
  wire[16:0] T3828;
  wire[16:0] T6932;
  wire[6:0] T3829;
  wire[9:0] T6933;
  wire T6934;
  wire T3830;
  wire T3831;
  wire[16:0] T3832;
  wire[16:0] T6935;
  wire[5:0] T3833;
  wire[5:0] T3834;
  wire[5:0] T6936;
  wire T3835;
  wire T3836;
  wire[10:0] T6937;
  wire T6938;
  wire[16:0] T3837;
  wire[16:0] T6939;
  wire[5:0] T3838;
  wire[10:0] T6940;
  wire T6941;
  wire T3839;
  wire T3840;
  wire[16:0] T3841;
  wire[16:0] T6942;
  wire[4:0] T3842;
  wire[4:0] T3843;
  wire[4:0] T6943;
  wire T3844;
  wire T3845;
  wire[11:0] T6944;
  wire T6945;
  wire[16:0] T3846;
  wire[16:0] T6946;
  wire[4:0] T3847;
  wire[11:0] T6947;
  wire T6948;
  wire T3848;
  wire T3849;
  wire[16:0] T3850;
  wire[16:0] T6949;
  wire[3:0] T3851;
  wire[3:0] T3852;
  wire[3:0] T6950;
  wire T3853;
  wire T3854;
  wire[12:0] T6951;
  wire T6952;
  wire[16:0] T3855;
  wire[16:0] T6953;
  wire[3:0] T3856;
  wire[12:0] T6954;
  wire T6955;
  wire T3857;
  wire T3858;
  wire[16:0] T3859;
  wire[16:0] T6956;
  wire[2:0] T3860;
  wire[2:0] T3861;
  wire[2:0] T6957;
  wire T3862;
  wire T3863;
  wire[13:0] T6958;
  wire T6959;
  wire[16:0] T3864;
  wire[16:0] T6960;
  wire[2:0] T3865;
  wire[13:0] T6961;
  wire T6962;
  wire T3866;
  wire T3867;
  wire[16:0] T3868;
  wire[16:0] T6963;
  wire[1:0] T3869;
  wire[1:0] T3870;
  wire[1:0] T6964;
  wire T3871;
  wire T3872;
  wire[14:0] T6965;
  wire T6966;
  wire[16:0] T3873;
  wire[16:0] T6967;
  wire[1:0] T3874;
  wire[14:0] T6968;
  wire T6969;
  wire T3875;
  wire T3876;
  wire[15:0] V_wire_en_16;
  wire[15:0] T6970;
  wire[16:0] T3877;
  wire[16:0] T3878;
  wire[16:0] T3879;
  wire[16:0] T3880;
  wire[16:0] T3881;
  wire[16:0] T3882;
  wire[16:0] T3883;
  wire[16:0] T3884;
  wire[16:0] T3885;
  wire[16:0] T3886;
  wire[16:0] T3887;
  wire[16:0] T3888;
  wire[16:0] T3889;
  wire[16:0] T3890;
  wire[16:0] T3891;
  wire[16:0] T3892;
  wire[16:0] T3893;
  wire[16:0] T3894;
  wire[16:0] T3895;
  wire[16:0] T6971;
  wire T3896;
  wire T3897;
  wire[16:0] T3898;
  wire[16:0] T3899;
  wire T3900;
  wire T3901;
  wire[3:0] T3902;
  wire T3903;
  wire T3904;
  wire[16:0] T3905;
  wire[16:0] T6972;
  wire[15:0] T3906;
  wire[15:0] T3907;
  wire[15:0] T6973;
  wire T3908;
  wire T3909;
  wire T6974;
  wire[16:0] T3910;
  wire[16:0] T6975;
  wire[15:0] T3911;
  wire T6976;
  wire T3912;
  wire T3913;
  wire[16:0] T3914;
  wire[16:0] T6977;
  wire[14:0] T3915;
  wire[14:0] T3916;
  wire[14:0] T6978;
  wire T3917;
  wire T3918;
  wire[1:0] T6979;
  wire T6980;
  wire[16:0] T3919;
  wire[16:0] T6981;
  wire[14:0] T3920;
  wire[1:0] T6982;
  wire T6983;
  wire T3921;
  wire T3922;
  wire[16:0] T3923;
  wire[16:0] T6984;
  wire[13:0] T3924;
  wire[13:0] T3925;
  wire[13:0] T6985;
  wire T3926;
  wire T3927;
  wire[2:0] T6986;
  wire T6987;
  wire[16:0] T3928;
  wire[16:0] T6988;
  wire[13:0] T3929;
  wire[2:0] T6989;
  wire T6990;
  wire T3930;
  wire T3931;
  wire[16:0] T3932;
  wire[16:0] T6991;
  wire[12:0] T3933;
  wire[12:0] T3934;
  wire[12:0] T6992;
  wire T3935;
  wire T3936;
  wire[3:0] T6993;
  wire T6994;
  wire[16:0] T3937;
  wire[16:0] T6995;
  wire[12:0] T3938;
  wire[3:0] T6996;
  wire T6997;
  wire T3939;
  wire T3940;
  wire[16:0] T3941;
  wire[16:0] T6998;
  wire[11:0] T3942;
  wire[11:0] T3943;
  wire[11:0] T6999;
  wire T3944;
  wire T3945;
  wire[4:0] T7000;
  wire T7001;
  wire[16:0] T3946;
  wire[16:0] T7002;
  wire[11:0] T3947;
  wire[4:0] T7003;
  wire T7004;
  wire T3948;
  wire T3949;
  wire[16:0] T3950;
  wire[16:0] T7005;
  wire[10:0] T3951;
  wire[10:0] T3952;
  wire[10:0] T7006;
  wire T3953;
  wire T3954;
  wire[5:0] T7007;
  wire T7008;
  wire[16:0] T3955;
  wire[16:0] T7009;
  wire[10:0] T3956;
  wire[5:0] T7010;
  wire T7011;
  wire T3957;
  wire T3958;
  wire[16:0] T3959;
  wire[16:0] T7012;
  wire[9:0] T3960;
  wire[9:0] T3961;
  wire[9:0] T7013;
  wire T3962;
  wire T3963;
  wire[6:0] T7014;
  wire T7015;
  wire[16:0] T3964;
  wire[16:0] T7016;
  wire[9:0] T3965;
  wire[6:0] T7017;
  wire T7018;
  wire T3966;
  wire T3967;
  wire[16:0] T3968;
  wire[16:0] T7019;
  wire[8:0] T3969;
  wire[8:0] T3970;
  wire[8:0] T7020;
  wire T3971;
  wire T3972;
  wire[7:0] T7021;
  wire T7022;
  wire[16:0] T3973;
  wire[16:0] T7023;
  wire[8:0] T3974;
  wire[7:0] T7024;
  wire T7025;
  wire T3975;
  wire T3976;
  wire[16:0] T3977;
  wire[16:0] T7026;
  wire[7:0] T3978;
  wire[7:0] T3979;
  wire[7:0] T7027;
  wire T3980;
  wire T3981;
  wire[8:0] T7028;
  wire T7029;
  wire[16:0] T3982;
  wire[16:0] T7030;
  wire[7:0] T3983;
  wire[8:0] T7031;
  wire T7032;
  wire T3984;
  wire T3985;
  wire[16:0] T3986;
  wire[16:0] T7033;
  wire[6:0] T3987;
  wire[6:0] T3988;
  wire[6:0] T7034;
  wire T3989;
  wire T3990;
  wire[9:0] T7035;
  wire T7036;
  wire[16:0] T3991;
  wire[16:0] T7037;
  wire[6:0] T3992;
  wire[9:0] T7038;
  wire T7039;
  wire T3993;
  wire T3994;
  wire[16:0] T3995;
  wire[16:0] T7040;
  wire[5:0] T3996;
  wire[5:0] T3997;
  wire[5:0] T7041;
  wire T3998;
  wire T3999;
  wire[10:0] T7042;
  wire T7043;
  wire[16:0] T4000;
  wire[16:0] T7044;
  wire[5:0] T4001;
  wire[10:0] T7045;
  wire T7046;
  wire T4002;
  wire T4003;
  wire[16:0] T4004;
  wire[16:0] T7047;
  wire[4:0] T4005;
  wire[4:0] T4006;
  wire[4:0] T7048;
  wire T4007;
  wire T4008;
  wire[11:0] T7049;
  wire T7050;
  wire[16:0] T4009;
  wire[16:0] T7051;
  wire[4:0] T4010;
  wire[11:0] T7052;
  wire T7053;
  wire T4011;
  wire T4012;
  wire[16:0] T4013;
  wire[16:0] T7054;
  wire[3:0] T4014;
  wire[3:0] T4015;
  wire[3:0] T7055;
  wire T4016;
  wire T4017;
  wire[12:0] T7056;
  wire T7057;
  wire[16:0] T4018;
  wire[16:0] T7058;
  wire[3:0] T4019;
  wire[12:0] T7059;
  wire T7060;
  wire T4020;
  wire T4021;
  wire[16:0] T4022;
  wire[16:0] T7061;
  wire[2:0] T4023;
  wire[2:0] T4024;
  wire[2:0] T7062;
  wire T4025;
  wire T4026;
  wire[13:0] T7063;
  wire T7064;
  wire[16:0] T4027;
  wire[16:0] T7065;
  wire[2:0] T4028;
  wire[13:0] T7066;
  wire T7067;
  wire T4029;
  wire T4030;
  wire[16:0] T4031;
  wire[16:0] T7068;
  wire[1:0] T4032;
  wire[1:0] T4033;
  wire[1:0] T7069;
  wire T4034;
  wire T4035;
  wire[14:0] T7070;
  wire T7071;
  wire[16:0] T4036;
  wire[16:0] T7072;
  wire[1:0] T4037;
  wire[14:0] T7073;
  wire T7074;
  wire T4038;
  wire T4039;
  wire[15:0] V_wire_en_17;
  wire[15:0] T7075;
  wire[16:0] T4040;
  wire[16:0] T4041;
  wire[16:0] T4042;
  wire[16:0] T4043;
  wire[16:0] T4044;
  wire[16:0] T4045;
  wire[16:0] T4046;
  wire[16:0] T4047;
  wire[16:0] T4048;
  wire[16:0] T4049;
  wire[16:0] T4050;
  wire[16:0] T4051;
  wire[16:0] T4052;
  wire[16:0] T4053;
  wire[16:0] T4054;
  wire[16:0] T4055;
  wire[16:0] T4056;
  wire[16:0] T4057;
  wire[16:0] T4058;
  wire[16:0] T7076;
  wire T4059;
  wire T4060;
  wire[16:0] T4061;
  wire[16:0] T4062;
  wire T4063;
  wire T4064;
  wire[3:0] T4065;
  wire T4066;
  wire T4067;
  wire[16:0] T4068;
  wire[16:0] T7077;
  wire[15:0] T4069;
  wire[15:0] T4070;
  wire[15:0] T7078;
  wire T4071;
  wire T4072;
  wire T7079;
  wire[16:0] T4073;
  wire[16:0] T7080;
  wire[15:0] T4074;
  wire T7081;
  wire T4075;
  wire T4076;
  wire[16:0] T4077;
  wire[16:0] T7082;
  wire[14:0] T4078;
  wire[14:0] T4079;
  wire[14:0] T7083;
  wire T4080;
  wire T4081;
  wire[1:0] T7084;
  wire T7085;
  wire[16:0] T4082;
  wire[16:0] T7086;
  wire[14:0] T4083;
  wire[1:0] T7087;
  wire T7088;
  wire T4084;
  wire T4085;
  wire[16:0] T4086;
  wire[16:0] T7089;
  wire[13:0] T4087;
  wire[13:0] T4088;
  wire[13:0] T7090;
  wire T4089;
  wire T4090;
  wire[2:0] T7091;
  wire T7092;
  wire[16:0] T4091;
  wire[16:0] T7093;
  wire[13:0] T4092;
  wire[2:0] T7094;
  wire T7095;
  wire T4093;
  wire T4094;
  wire[16:0] T4095;
  wire[16:0] T7096;
  wire[12:0] T4096;
  wire[12:0] T4097;
  wire[12:0] T7097;
  wire T4098;
  wire T4099;
  wire[3:0] T7098;
  wire T7099;
  wire[16:0] T4100;
  wire[16:0] T7100;
  wire[12:0] T4101;
  wire[3:0] T7101;
  wire T7102;
  wire T4102;
  wire T4103;
  wire[16:0] T4104;
  wire[16:0] T7103;
  wire[11:0] T4105;
  wire[11:0] T4106;
  wire[11:0] T7104;
  wire T4107;
  wire T4108;
  wire[4:0] T7105;
  wire T7106;
  wire[16:0] T4109;
  wire[16:0] T7107;
  wire[11:0] T4110;
  wire[4:0] T7108;
  wire T7109;
  wire T4111;
  wire T4112;
  wire[16:0] T4113;
  wire[16:0] T7110;
  wire[10:0] T4114;
  wire[10:0] T4115;
  wire[10:0] T7111;
  wire T4116;
  wire T4117;
  wire[5:0] T7112;
  wire T7113;
  wire[16:0] T4118;
  wire[16:0] T7114;
  wire[10:0] T4119;
  wire[5:0] T7115;
  wire T7116;
  wire T4120;
  wire T4121;
  wire[16:0] T4122;
  wire[16:0] T7117;
  wire[9:0] T4123;
  wire[9:0] T4124;
  wire[9:0] T7118;
  wire T4125;
  wire T4126;
  wire[6:0] T7119;
  wire T7120;
  wire[16:0] T4127;
  wire[16:0] T7121;
  wire[9:0] T4128;
  wire[6:0] T7122;
  wire T7123;
  wire T4129;
  wire T4130;
  wire[16:0] T4131;
  wire[16:0] T7124;
  wire[8:0] T4132;
  wire[8:0] T4133;
  wire[8:0] T7125;
  wire T4134;
  wire T4135;
  wire[7:0] T7126;
  wire T7127;
  wire[16:0] T4136;
  wire[16:0] T7128;
  wire[8:0] T4137;
  wire[7:0] T7129;
  wire T7130;
  wire T4138;
  wire T4139;
  wire[16:0] T4140;
  wire[16:0] T7131;
  wire[7:0] T4141;
  wire[7:0] T4142;
  wire[7:0] T7132;
  wire T4143;
  wire T4144;
  wire[8:0] T7133;
  wire T7134;
  wire[16:0] T4145;
  wire[16:0] T7135;
  wire[7:0] T4146;
  wire[8:0] T7136;
  wire T7137;
  wire T4147;
  wire T4148;
  wire[16:0] T4149;
  wire[16:0] T7138;
  wire[6:0] T4150;
  wire[6:0] T4151;
  wire[6:0] T7139;
  wire T4152;
  wire T4153;
  wire[9:0] T7140;
  wire T7141;
  wire[16:0] T4154;
  wire[16:0] T7142;
  wire[6:0] T4155;
  wire[9:0] T7143;
  wire T7144;
  wire T4156;
  wire T4157;
  wire[16:0] T4158;
  wire[16:0] T7145;
  wire[5:0] T4159;
  wire[5:0] T4160;
  wire[5:0] T7146;
  wire T4161;
  wire T4162;
  wire[10:0] T7147;
  wire T7148;
  wire[16:0] T4163;
  wire[16:0] T7149;
  wire[5:0] T4164;
  wire[10:0] T7150;
  wire T7151;
  wire T4165;
  wire T4166;
  wire[16:0] T4167;
  wire[16:0] T7152;
  wire[4:0] T4168;
  wire[4:0] T4169;
  wire[4:0] T7153;
  wire T4170;
  wire T4171;
  wire[11:0] T7154;
  wire T7155;
  wire[16:0] T4172;
  wire[16:0] T7156;
  wire[4:0] T4173;
  wire[11:0] T7157;
  wire T7158;
  wire T4174;
  wire T4175;
  wire[16:0] T4176;
  wire[16:0] T7159;
  wire[3:0] T4177;
  wire[3:0] T4178;
  wire[3:0] T7160;
  wire T4179;
  wire T4180;
  wire[12:0] T7161;
  wire T7162;
  wire[16:0] T4181;
  wire[16:0] T7163;
  wire[3:0] T4182;
  wire[12:0] T7164;
  wire T7165;
  wire T4183;
  wire T4184;
  wire[16:0] T4185;
  wire[16:0] T7166;
  wire[2:0] T4186;
  wire[2:0] T4187;
  wire[2:0] T7167;
  wire T4188;
  wire T4189;
  wire[13:0] T7168;
  wire T7169;
  wire[16:0] T4190;
  wire[16:0] T7170;
  wire[2:0] T4191;
  wire[13:0] T7171;
  wire T7172;
  wire T4192;
  wire T4193;
  wire[16:0] T4194;
  wire[16:0] T7173;
  wire[1:0] T4195;
  wire[1:0] T4196;
  wire[1:0] T7174;
  wire T4197;
  wire T4198;
  wire[14:0] T7175;
  wire T7176;
  wire[16:0] T4199;
  wire[16:0] T7177;
  wire[1:0] T4200;
  wire[14:0] T7178;
  wire T7179;
  wire T4201;
  wire T4202;
  wire[15:0] V_wire_en_18;
  wire[15:0] T7180;
  wire[16:0] T4203;
  wire[16:0] T4204;
  wire[16:0] T4205;
  wire[16:0] T4206;
  wire[16:0] T4207;
  wire[16:0] T4208;
  wire[16:0] T4209;
  wire[16:0] T4210;
  wire[16:0] T4211;
  wire[16:0] T4212;
  wire[16:0] T4213;
  wire[16:0] T4214;
  wire[16:0] T4215;
  wire[16:0] T4216;
  wire[16:0] T4217;
  wire[16:0] T4218;
  wire[16:0] T4219;
  wire[16:0] T4220;
  wire[16:0] T4221;
  wire[16:0] T7181;
  wire T4222;
  wire T4223;
  wire[16:0] T4224;
  wire[16:0] T4225;
  wire T4226;
  wire T4227;
  wire[3:0] T4228;
  wire T4229;
  wire T4230;
  wire[16:0] T4231;
  wire[16:0] T7182;
  wire[15:0] T4232;
  wire[15:0] T4233;
  wire[15:0] T7183;
  wire T4234;
  wire T4235;
  wire T7184;
  wire[16:0] T4236;
  wire[16:0] T7185;
  wire[15:0] T4237;
  wire T7186;
  wire T4238;
  wire T4239;
  wire[16:0] T4240;
  wire[16:0] T7187;
  wire[14:0] T4241;
  wire[14:0] T4242;
  wire[14:0] T7188;
  wire T4243;
  wire T4244;
  wire[1:0] T7189;
  wire T7190;
  wire[16:0] T4245;
  wire[16:0] T7191;
  wire[14:0] T4246;
  wire[1:0] T7192;
  wire T7193;
  wire T4247;
  wire T4248;
  wire[16:0] T4249;
  wire[16:0] T7194;
  wire[13:0] T4250;
  wire[13:0] T4251;
  wire[13:0] T7195;
  wire T4252;
  wire T4253;
  wire[2:0] T7196;
  wire T7197;
  wire[16:0] T4254;
  wire[16:0] T7198;
  wire[13:0] T4255;
  wire[2:0] T7199;
  wire T7200;
  wire T4256;
  wire T4257;
  wire[16:0] T4258;
  wire[16:0] T7201;
  wire[12:0] T4259;
  wire[12:0] T4260;
  wire[12:0] T7202;
  wire T4261;
  wire T4262;
  wire[3:0] T7203;
  wire T7204;
  wire[16:0] T4263;
  wire[16:0] T7205;
  wire[12:0] T4264;
  wire[3:0] T7206;
  wire T7207;
  wire T4265;
  wire T4266;
  wire[16:0] T4267;
  wire[16:0] T7208;
  wire[11:0] T4268;
  wire[11:0] T4269;
  wire[11:0] T7209;
  wire T4270;
  wire T4271;
  wire[4:0] T7210;
  wire T7211;
  wire[16:0] T4272;
  wire[16:0] T7212;
  wire[11:0] T4273;
  wire[4:0] T7213;
  wire T7214;
  wire T4274;
  wire T4275;
  wire[16:0] T4276;
  wire[16:0] T7215;
  wire[10:0] T4277;
  wire[10:0] T4278;
  wire[10:0] T7216;
  wire T4279;
  wire T4280;
  wire[5:0] T7217;
  wire T7218;
  wire[16:0] T4281;
  wire[16:0] T7219;
  wire[10:0] T4282;
  wire[5:0] T7220;
  wire T7221;
  wire T4283;
  wire T4284;
  wire[16:0] T4285;
  wire[16:0] T7222;
  wire[9:0] T4286;
  wire[9:0] T4287;
  wire[9:0] T7223;
  wire T4288;
  wire T4289;
  wire[6:0] T7224;
  wire T7225;
  wire[16:0] T4290;
  wire[16:0] T7226;
  wire[9:0] T4291;
  wire[6:0] T7227;
  wire T7228;
  wire T4292;
  wire T4293;
  wire[16:0] T4294;
  wire[16:0] T7229;
  wire[8:0] T4295;
  wire[8:0] T4296;
  wire[8:0] T7230;
  wire T4297;
  wire T4298;
  wire[7:0] T7231;
  wire T7232;
  wire[16:0] T4299;
  wire[16:0] T7233;
  wire[8:0] T4300;
  wire[7:0] T7234;
  wire T7235;
  wire T4301;
  wire T4302;
  wire[16:0] T4303;
  wire[16:0] T7236;
  wire[7:0] T4304;
  wire[7:0] T4305;
  wire[7:0] T7237;
  wire T4306;
  wire T4307;
  wire[8:0] T7238;
  wire T7239;
  wire[16:0] T4308;
  wire[16:0] T7240;
  wire[7:0] T4309;
  wire[8:0] T7241;
  wire T7242;
  wire T4310;
  wire T4311;
  wire[16:0] T4312;
  wire[16:0] T7243;
  wire[6:0] T4313;
  wire[6:0] T4314;
  wire[6:0] T7244;
  wire T4315;
  wire T4316;
  wire[9:0] T7245;
  wire T7246;
  wire[16:0] T4317;
  wire[16:0] T7247;
  wire[6:0] T4318;
  wire[9:0] T7248;
  wire T7249;
  wire T4319;
  wire T4320;
  wire[16:0] T4321;
  wire[16:0] T7250;
  wire[5:0] T4322;
  wire[5:0] T4323;
  wire[5:0] T7251;
  wire T4324;
  wire T4325;
  wire[10:0] T7252;
  wire T7253;
  wire[16:0] T4326;
  wire[16:0] T7254;
  wire[5:0] T4327;
  wire[10:0] T7255;
  wire T7256;
  wire T4328;
  wire T4329;
  wire[16:0] T4330;
  wire[16:0] T7257;
  wire[4:0] T4331;
  wire[4:0] T4332;
  wire[4:0] T7258;
  wire T4333;
  wire T4334;
  wire[11:0] T7259;
  wire T7260;
  wire[16:0] T4335;
  wire[16:0] T7261;
  wire[4:0] T4336;
  wire[11:0] T7262;
  wire T7263;
  wire T4337;
  wire T4338;
  wire[16:0] T4339;
  wire[16:0] T7264;
  wire[3:0] T4340;
  wire[3:0] T4341;
  wire[3:0] T7265;
  wire T4342;
  wire T4343;
  wire[12:0] T7266;
  wire T7267;
  wire[16:0] T4344;
  wire[16:0] T7268;
  wire[3:0] T4345;
  wire[12:0] T7269;
  wire T7270;
  wire T4346;
  wire T4347;
  wire[16:0] T4348;
  wire[16:0] T7271;
  wire[2:0] T4349;
  wire[2:0] T4350;
  wire[2:0] T7272;
  wire T4351;
  wire T4352;
  wire[13:0] T7273;
  wire T7274;
  wire[16:0] T4353;
  wire[16:0] T7275;
  wire[2:0] T4354;
  wire[13:0] T7276;
  wire T7277;
  wire T4355;
  wire T4356;
  wire[16:0] T4357;
  wire[16:0] T7278;
  wire[1:0] T4358;
  wire[1:0] T4359;
  wire[1:0] T7279;
  wire T4360;
  wire T4361;
  wire[14:0] T7280;
  wire T7281;
  wire[16:0] T4362;
  wire[16:0] T7282;
  wire[1:0] T4363;
  wire[14:0] T7283;
  wire T7284;
  wire T4364;
  wire T4365;
  wire[15:0] V_wire_en_19;
  wire[15:0] T7285;
  wire[16:0] T4366;
  wire[16:0] T4367;
  wire[16:0] T4368;
  wire[16:0] T4369;
  wire[16:0] T4370;
  wire[16:0] T4371;
  wire[16:0] T4372;
  wire[16:0] T4373;
  wire[16:0] T4374;
  wire[16:0] T4375;
  wire[16:0] T4376;
  wire[16:0] T4377;
  wire[16:0] T4378;
  wire[16:0] T4379;
  wire[16:0] T4380;
  wire[16:0] T4381;
  wire[16:0] T4382;
  wire[16:0] T4383;
  wire[16:0] T4384;
  wire[16:0] T7286;
  wire T4385;
  wire T4386;
  wire[16:0] T4387;
  wire[16:0] T4388;
  wire T4389;
  wire T4390;
  wire[3:0] T4391;
  wire T4392;
  wire T4393;
  wire[16:0] T4394;
  wire[16:0] T7287;
  wire[15:0] T4395;
  wire[15:0] T4396;
  wire[15:0] T7288;
  wire T4397;
  wire T4398;
  wire T7289;
  wire[16:0] T4399;
  wire[16:0] T7290;
  wire[15:0] T4400;
  wire T7291;
  wire T4401;
  wire T4402;
  wire[16:0] T4403;
  wire[16:0] T7292;
  wire[14:0] T4404;
  wire[14:0] T4405;
  wire[14:0] T7293;
  wire T4406;
  wire T4407;
  wire[1:0] T7294;
  wire T7295;
  wire[16:0] T4408;
  wire[16:0] T7296;
  wire[14:0] T4409;
  wire[1:0] T7297;
  wire T7298;
  wire T4410;
  wire T4411;
  wire[16:0] T4412;
  wire[16:0] T7299;
  wire[13:0] T4413;
  wire[13:0] T4414;
  wire[13:0] T7300;
  wire T4415;
  wire T4416;
  wire[2:0] T7301;
  wire T7302;
  wire[16:0] T4417;
  wire[16:0] T7303;
  wire[13:0] T4418;
  wire[2:0] T7304;
  wire T7305;
  wire T4419;
  wire T4420;
  wire[16:0] T4421;
  wire[16:0] T7306;
  wire[12:0] T4422;
  wire[12:0] T4423;
  wire[12:0] T7307;
  wire T4424;
  wire T4425;
  wire[3:0] T7308;
  wire T7309;
  wire[16:0] T4426;
  wire[16:0] T7310;
  wire[12:0] T4427;
  wire[3:0] T7311;
  wire T7312;
  wire T4428;
  wire T4429;
  wire[16:0] T4430;
  wire[16:0] T7313;
  wire[11:0] T4431;
  wire[11:0] T4432;
  wire[11:0] T7314;
  wire T4433;
  wire T4434;
  wire[4:0] T7315;
  wire T7316;
  wire[16:0] T4435;
  wire[16:0] T7317;
  wire[11:0] T4436;
  wire[4:0] T7318;
  wire T7319;
  wire T4437;
  wire T4438;
  wire[16:0] T4439;
  wire[16:0] T7320;
  wire[10:0] T4440;
  wire[10:0] T4441;
  wire[10:0] T7321;
  wire T4442;
  wire T4443;
  wire[5:0] T7322;
  wire T7323;
  wire[16:0] T4444;
  wire[16:0] T7324;
  wire[10:0] T4445;
  wire[5:0] T7325;
  wire T7326;
  wire T4446;
  wire T4447;
  wire[16:0] T4448;
  wire[16:0] T7327;
  wire[9:0] T4449;
  wire[9:0] T4450;
  wire[9:0] T7328;
  wire T4451;
  wire T4452;
  wire[6:0] T7329;
  wire T7330;
  wire[16:0] T4453;
  wire[16:0] T7331;
  wire[9:0] T4454;
  wire[6:0] T7332;
  wire T7333;
  wire T4455;
  wire T4456;
  wire[16:0] T4457;
  wire[16:0] T7334;
  wire[8:0] T4458;
  wire[8:0] T4459;
  wire[8:0] T7335;
  wire T4460;
  wire T4461;
  wire[7:0] T7336;
  wire T7337;
  wire[16:0] T4462;
  wire[16:0] T7338;
  wire[8:0] T4463;
  wire[7:0] T7339;
  wire T7340;
  wire T4464;
  wire T4465;
  wire[16:0] T4466;
  wire[16:0] T7341;
  wire[7:0] T4467;
  wire[7:0] T4468;
  wire[7:0] T7342;
  wire T4469;
  wire T4470;
  wire[8:0] T7343;
  wire T7344;
  wire[16:0] T4471;
  wire[16:0] T7345;
  wire[7:0] T4472;
  wire[8:0] T7346;
  wire T7347;
  wire T4473;
  wire T4474;
  wire[16:0] T4475;
  wire[16:0] T7348;
  wire[6:0] T4476;
  wire[6:0] T4477;
  wire[6:0] T7349;
  wire T4478;
  wire T4479;
  wire[9:0] T7350;
  wire T7351;
  wire[16:0] T4480;
  wire[16:0] T7352;
  wire[6:0] T4481;
  wire[9:0] T7353;
  wire T7354;
  wire T4482;
  wire T4483;
  wire[16:0] T4484;
  wire[16:0] T7355;
  wire[5:0] T4485;
  wire[5:0] T4486;
  wire[5:0] T7356;
  wire T4487;
  wire T4488;
  wire[10:0] T7357;
  wire T7358;
  wire[16:0] T4489;
  wire[16:0] T7359;
  wire[5:0] T4490;
  wire[10:0] T7360;
  wire T7361;
  wire T4491;
  wire T4492;
  wire[16:0] T4493;
  wire[16:0] T7362;
  wire[4:0] T4494;
  wire[4:0] T4495;
  wire[4:0] T7363;
  wire T4496;
  wire T4497;
  wire[11:0] T7364;
  wire T7365;
  wire[16:0] T4498;
  wire[16:0] T7366;
  wire[4:0] T4499;
  wire[11:0] T7367;
  wire T7368;
  wire T4500;
  wire T4501;
  wire[16:0] T4502;
  wire[16:0] T7369;
  wire[3:0] T4503;
  wire[3:0] T4504;
  wire[3:0] T7370;
  wire T4505;
  wire T4506;
  wire[12:0] T7371;
  wire T7372;
  wire[16:0] T4507;
  wire[16:0] T7373;
  wire[3:0] T4508;
  wire[12:0] T7374;
  wire T7375;
  wire T4509;
  wire T4510;
  wire[16:0] T4511;
  wire[16:0] T7376;
  wire[2:0] T4512;
  wire[2:0] T4513;
  wire[2:0] T7377;
  wire T4514;
  wire T4515;
  wire[13:0] T7378;
  wire T7379;
  wire[16:0] T4516;
  wire[16:0] T7380;
  wire[2:0] T4517;
  wire[13:0] T7381;
  wire T7382;
  wire T4518;
  wire T4519;
  wire[16:0] T4520;
  wire[16:0] T7383;
  wire[1:0] T4521;
  wire[1:0] T4522;
  wire[1:0] T7384;
  wire T4523;
  wire T4524;
  wire[14:0] T7385;
  wire T7386;
  wire[16:0] T4525;
  wire[16:0] T7387;
  wire[1:0] T4526;
  wire[14:0] T7388;
  wire T7389;
  wire T4527;
  wire T4528;
  wire[15:0] V_wire_en_20;
  wire[15:0] T7390;
  wire[16:0] T4529;
  wire[16:0] T4530;
  wire[16:0] T4531;
  wire[16:0] T4532;
  wire[16:0] T4533;
  wire[16:0] T4534;
  wire[16:0] T4535;
  wire[16:0] T4536;
  wire[16:0] T4537;
  wire[16:0] T4538;
  wire[16:0] T4539;
  wire[16:0] T4540;
  wire[16:0] T4541;
  wire[16:0] T4542;
  wire[16:0] T4543;
  wire[16:0] T4544;
  wire[16:0] T4545;
  wire[16:0] T4546;
  wire[16:0] T4547;
  wire[16:0] T7391;
  wire T4548;
  wire T4549;
  wire[16:0] T4550;
  wire[16:0] T4551;
  wire T4552;
  wire T4553;
  wire[3:0] T4554;
  wire T4555;
  wire T4556;
  wire[16:0] T4557;
  wire[16:0] T7392;
  wire[15:0] T4558;
  wire[15:0] T4559;
  wire[15:0] T7393;
  wire T4560;
  wire T4561;
  wire T7394;
  wire[16:0] T4562;
  wire[16:0] T7395;
  wire[15:0] T4563;
  wire T7396;
  wire T4564;
  wire T4565;
  wire[16:0] T4566;
  wire[16:0] T7397;
  wire[14:0] T4567;
  wire[14:0] T4568;
  wire[14:0] T7398;
  wire T4569;
  wire T4570;
  wire[1:0] T7399;
  wire T7400;
  wire[16:0] T4571;
  wire[16:0] T7401;
  wire[14:0] T4572;
  wire[1:0] T7402;
  wire T7403;
  wire T4573;
  wire T4574;
  wire[16:0] T4575;
  wire[16:0] T7404;
  wire[13:0] T4576;
  wire[13:0] T4577;
  wire[13:0] T7405;
  wire T4578;
  wire T4579;
  wire[2:0] T7406;
  wire T7407;
  wire[16:0] T4580;
  wire[16:0] T7408;
  wire[13:0] T4581;
  wire[2:0] T7409;
  wire T7410;
  wire T4582;
  wire T4583;
  wire[16:0] T4584;
  wire[16:0] T7411;
  wire[12:0] T4585;
  wire[12:0] T4586;
  wire[12:0] T7412;
  wire T4587;
  wire T4588;
  wire[3:0] T7413;
  wire T7414;
  wire[16:0] T4589;
  wire[16:0] T7415;
  wire[12:0] T4590;
  wire[3:0] T7416;
  wire T7417;
  wire T4591;
  wire T4592;
  wire[16:0] T4593;
  wire[16:0] T7418;
  wire[11:0] T4594;
  wire[11:0] T4595;
  wire[11:0] T7419;
  wire T4596;
  wire T4597;
  wire[4:0] T7420;
  wire T7421;
  wire[16:0] T4598;
  wire[16:0] T7422;
  wire[11:0] T4599;
  wire[4:0] T7423;
  wire T7424;
  wire T4600;
  wire T4601;
  wire[16:0] T4602;
  wire[16:0] T7425;
  wire[10:0] T4603;
  wire[10:0] T4604;
  wire[10:0] T7426;
  wire T4605;
  wire T4606;
  wire[5:0] T7427;
  wire T7428;
  wire[16:0] T4607;
  wire[16:0] T7429;
  wire[10:0] T4608;
  wire[5:0] T7430;
  wire T7431;
  wire T4609;
  wire T4610;
  wire[16:0] T4611;
  wire[16:0] T7432;
  wire[9:0] T4612;
  wire[9:0] T4613;
  wire[9:0] T7433;
  wire T4614;
  wire T4615;
  wire[6:0] T7434;
  wire T7435;
  wire[16:0] T4616;
  wire[16:0] T7436;
  wire[9:0] T4617;
  wire[6:0] T7437;
  wire T7438;
  wire T4618;
  wire T4619;
  wire[16:0] T4620;
  wire[16:0] T7439;
  wire[8:0] T4621;
  wire[8:0] T4622;
  wire[8:0] T7440;
  wire T4623;
  wire T4624;
  wire[7:0] T7441;
  wire T7442;
  wire[16:0] T4625;
  wire[16:0] T7443;
  wire[8:0] T4626;
  wire[7:0] T7444;
  wire T7445;
  wire T4627;
  wire T4628;
  wire[16:0] T4629;
  wire[16:0] T7446;
  wire[7:0] T4630;
  wire[7:0] T4631;
  wire[7:0] T7447;
  wire T4632;
  wire T4633;
  wire[8:0] T7448;
  wire T7449;
  wire[16:0] T4634;
  wire[16:0] T7450;
  wire[7:0] T4635;
  wire[8:0] T7451;
  wire T7452;
  wire T4636;
  wire T4637;
  wire[16:0] T4638;
  wire[16:0] T7453;
  wire[6:0] T4639;
  wire[6:0] T4640;
  wire[6:0] T7454;
  wire T4641;
  wire T4642;
  wire[9:0] T7455;
  wire T7456;
  wire[16:0] T4643;
  wire[16:0] T7457;
  wire[6:0] T4644;
  wire[9:0] T7458;
  wire T7459;
  wire T4645;
  wire T4646;
  wire[16:0] T4647;
  wire[16:0] T7460;
  wire[5:0] T4648;
  wire[5:0] T4649;
  wire[5:0] T7461;
  wire T4650;
  wire T4651;
  wire[10:0] T7462;
  wire T7463;
  wire[16:0] T4652;
  wire[16:0] T7464;
  wire[5:0] T4653;
  wire[10:0] T7465;
  wire T7466;
  wire T4654;
  wire T4655;
  wire[16:0] T4656;
  wire[16:0] T7467;
  wire[4:0] T4657;
  wire[4:0] T4658;
  wire[4:0] T7468;
  wire T4659;
  wire T4660;
  wire[11:0] T7469;
  wire T7470;
  wire[16:0] T4661;
  wire[16:0] T7471;
  wire[4:0] T4662;
  wire[11:0] T7472;
  wire T7473;
  wire T4663;
  wire T4664;
  wire[16:0] T4665;
  wire[16:0] T7474;
  wire[3:0] T4666;
  wire[3:0] T4667;
  wire[3:0] T7475;
  wire T4668;
  wire T4669;
  wire[12:0] T7476;
  wire T7477;
  wire[16:0] T4670;
  wire[16:0] T7478;
  wire[3:0] T4671;
  wire[12:0] T7479;
  wire T7480;
  wire T4672;
  wire T4673;
  wire[16:0] T4674;
  wire[16:0] T7481;
  wire[2:0] T4675;
  wire[2:0] T4676;
  wire[2:0] T7482;
  wire T4677;
  wire T4678;
  wire[13:0] T7483;
  wire T7484;
  wire[16:0] T4679;
  wire[16:0] T7485;
  wire[2:0] T4680;
  wire[13:0] T7486;
  wire T7487;
  wire T4681;
  wire T4682;
  wire[16:0] T4683;
  wire[16:0] T7488;
  wire[1:0] T4684;
  wire[1:0] T4685;
  wire[1:0] T7489;
  wire T4686;
  wire T4687;
  wire[14:0] T7490;
  wire T7491;
  wire[16:0] T4688;
  wire[16:0] T7492;
  wire[1:0] T4689;
  wire[14:0] T7493;
  wire T7494;
  wire T4690;
  wire T4691;
  wire[15:0] V_wire_en_21;
  wire[15:0] T7495;
  wire[16:0] T4692;
  wire[16:0] T4693;
  wire[16:0] T4694;
  wire[16:0] T4695;
  wire[16:0] T4696;
  wire[16:0] T4697;
  wire[16:0] T4698;
  wire[16:0] T4699;
  wire[16:0] T4700;
  wire[16:0] T4701;
  wire[16:0] T4702;
  wire[16:0] T4703;
  wire[16:0] T4704;
  wire[16:0] T4705;
  wire[16:0] T4706;
  wire[16:0] T4707;
  wire[16:0] T4708;
  wire[16:0] T4709;
  wire[16:0] T4710;
  wire[16:0] T7496;
  wire T4711;
  wire T4712;
  wire[16:0] T4713;
  wire[16:0] T4714;
  wire T4715;
  wire T4716;
  wire[3:0] T4717;
  wire T4718;
  wire T4719;
  wire[16:0] T4720;
  wire[16:0] T7497;
  wire[15:0] T4721;
  wire[15:0] T4722;
  wire[15:0] T7498;
  wire T4723;
  wire T4724;
  wire T7499;
  wire[16:0] T4725;
  wire[16:0] T7500;
  wire[15:0] T4726;
  wire T7501;
  wire T4727;
  wire T4728;
  wire[16:0] T4729;
  wire[16:0] T7502;
  wire[14:0] T4730;
  wire[14:0] T4731;
  wire[14:0] T7503;
  wire T4732;
  wire T4733;
  wire[1:0] T7504;
  wire T7505;
  wire[16:0] T4734;
  wire[16:0] T7506;
  wire[14:0] T4735;
  wire[1:0] T7507;
  wire T7508;
  wire T4736;
  wire T4737;
  wire[16:0] T4738;
  wire[16:0] T7509;
  wire[13:0] T4739;
  wire[13:0] T4740;
  wire[13:0] T7510;
  wire T4741;
  wire T4742;
  wire[2:0] T7511;
  wire T7512;
  wire[16:0] T4743;
  wire[16:0] T7513;
  wire[13:0] T4744;
  wire[2:0] T7514;
  wire T7515;
  wire T4745;
  wire T4746;
  wire[16:0] T4747;
  wire[16:0] T7516;
  wire[12:0] T4748;
  wire[12:0] T4749;
  wire[12:0] T7517;
  wire T4750;
  wire T4751;
  wire[3:0] T7518;
  wire T7519;
  wire[16:0] T4752;
  wire[16:0] T7520;
  wire[12:0] T4753;
  wire[3:0] T7521;
  wire T7522;
  wire T4754;
  wire T4755;
  wire[16:0] T4756;
  wire[16:0] T7523;
  wire[11:0] T4757;
  wire[11:0] T4758;
  wire[11:0] T7524;
  wire T4759;
  wire T4760;
  wire[4:0] T7525;
  wire T7526;
  wire[16:0] T4761;
  wire[16:0] T7527;
  wire[11:0] T4762;
  wire[4:0] T7528;
  wire T7529;
  wire T4763;
  wire T4764;
  wire[16:0] T4765;
  wire[16:0] T7530;
  wire[10:0] T4766;
  wire[10:0] T4767;
  wire[10:0] T7531;
  wire T4768;
  wire T4769;
  wire[5:0] T7532;
  wire T7533;
  wire[16:0] T4770;
  wire[16:0] T7534;
  wire[10:0] T4771;
  wire[5:0] T7535;
  wire T7536;
  wire T4772;
  wire T4773;
  wire[16:0] T4774;
  wire[16:0] T7537;
  wire[9:0] T4775;
  wire[9:0] T4776;
  wire[9:0] T7538;
  wire T4777;
  wire T4778;
  wire[6:0] T7539;
  wire T7540;
  wire[16:0] T4779;
  wire[16:0] T7541;
  wire[9:0] T4780;
  wire[6:0] T7542;
  wire T7543;
  wire T4781;
  wire T4782;
  wire[16:0] T4783;
  wire[16:0] T7544;
  wire[8:0] T4784;
  wire[8:0] T4785;
  wire[8:0] T7545;
  wire T4786;
  wire T4787;
  wire[7:0] T7546;
  wire T7547;
  wire[16:0] T4788;
  wire[16:0] T7548;
  wire[8:0] T4789;
  wire[7:0] T7549;
  wire T7550;
  wire T4790;
  wire T4791;
  wire[16:0] T4792;
  wire[16:0] T7551;
  wire[7:0] T4793;
  wire[7:0] T4794;
  wire[7:0] T7552;
  wire T4795;
  wire T4796;
  wire[8:0] T7553;
  wire T7554;
  wire[16:0] T4797;
  wire[16:0] T7555;
  wire[7:0] T4798;
  wire[8:0] T7556;
  wire T7557;
  wire T4799;
  wire T4800;
  wire[16:0] T4801;
  wire[16:0] T7558;
  wire[6:0] T4802;
  wire[6:0] T4803;
  wire[6:0] T7559;
  wire T4804;
  wire T4805;
  wire[9:0] T7560;
  wire T7561;
  wire[16:0] T4806;
  wire[16:0] T7562;
  wire[6:0] T4807;
  wire[9:0] T7563;
  wire T7564;
  wire T4808;
  wire T4809;
  wire[16:0] T4810;
  wire[16:0] T7565;
  wire[5:0] T4811;
  wire[5:0] T4812;
  wire[5:0] T7566;
  wire T4813;
  wire T4814;
  wire[10:0] T7567;
  wire T7568;
  wire[16:0] T4815;
  wire[16:0] T7569;
  wire[5:0] T4816;
  wire[10:0] T7570;
  wire T7571;
  wire T4817;
  wire T4818;
  wire[16:0] T4819;
  wire[16:0] T7572;
  wire[4:0] T4820;
  wire[4:0] T4821;
  wire[4:0] T7573;
  wire T4822;
  wire T4823;
  wire[11:0] T7574;
  wire T7575;
  wire[16:0] T4824;
  wire[16:0] T7576;
  wire[4:0] T4825;
  wire[11:0] T7577;
  wire T7578;
  wire T4826;
  wire T4827;
  wire[16:0] T4828;
  wire[16:0] T7579;
  wire[3:0] T4829;
  wire[3:0] T4830;
  wire[3:0] T7580;
  wire T4831;
  wire T4832;
  wire[12:0] T7581;
  wire T7582;
  wire[16:0] T4833;
  wire[16:0] T7583;
  wire[3:0] T4834;
  wire[12:0] T7584;
  wire T7585;
  wire T4835;
  wire T4836;
  wire[16:0] T4837;
  wire[16:0] T7586;
  wire[2:0] T4838;
  wire[2:0] T4839;
  wire[2:0] T7587;
  wire T4840;
  wire T4841;
  wire[13:0] T7588;
  wire T7589;
  wire[16:0] T4842;
  wire[16:0] T7590;
  wire[2:0] T4843;
  wire[13:0] T7591;
  wire T7592;
  wire T4844;
  wire T4845;
  wire[16:0] T4846;
  wire[16:0] T7593;
  wire[1:0] T4847;
  wire[1:0] T4848;
  wire[1:0] T7594;
  wire T4849;
  wire T4850;
  wire[14:0] T7595;
  wire T7596;
  wire[16:0] T4851;
  wire[16:0] T7597;
  wire[1:0] T4852;
  wire[14:0] T7598;
  wire T7599;
  wire T4853;
  wire T4854;
  wire[15:0] V_wire_en_22;
  wire[15:0] T7600;
  wire[16:0] T4855;
  wire[16:0] T4856;
  wire[16:0] T4857;
  wire[16:0] T4858;
  wire[16:0] T4859;
  wire[16:0] T4860;
  wire[16:0] T4861;
  wire[16:0] T4862;
  wire[16:0] T4863;
  wire[16:0] T4864;
  wire[16:0] T4865;
  wire[16:0] T4866;
  wire[16:0] T4867;
  wire[16:0] T4868;
  wire[16:0] T4869;
  wire[16:0] T4870;
  wire[16:0] T4871;
  wire[16:0] T4872;
  wire[16:0] T4873;
  wire[16:0] T7601;
  wire T4874;
  wire T4875;
  wire[16:0] T4876;
  wire[16:0] T4877;
  wire T4878;
  wire T4879;
  wire[3:0] T4880;
  wire T4881;
  wire T4882;
  wire[16:0] T4883;
  wire[16:0] T7602;
  wire[15:0] T4884;
  wire[15:0] T4885;
  wire[15:0] T7603;
  wire T4886;
  wire T4887;
  wire T7604;
  wire[16:0] T4888;
  wire[16:0] T7605;
  wire[15:0] T4889;
  wire T7606;
  wire T4890;
  wire T4891;
  wire[16:0] T4892;
  wire[16:0] T7607;
  wire[14:0] T4893;
  wire[14:0] T4894;
  wire[14:0] T7608;
  wire T4895;
  wire T4896;
  wire[1:0] T7609;
  wire T7610;
  wire[16:0] T4897;
  wire[16:0] T7611;
  wire[14:0] T4898;
  wire[1:0] T7612;
  wire T7613;
  wire T4899;
  wire T4900;
  wire[16:0] T4901;
  wire[16:0] T7614;
  wire[13:0] T4902;
  wire[13:0] T4903;
  wire[13:0] T7615;
  wire T4904;
  wire T4905;
  wire[2:0] T7616;
  wire T7617;
  wire[16:0] T4906;
  wire[16:0] T7618;
  wire[13:0] T4907;
  wire[2:0] T7619;
  wire T7620;
  wire T4908;
  wire T4909;
  wire[16:0] T4910;
  wire[16:0] T7621;
  wire[12:0] T4911;
  wire[12:0] T4912;
  wire[12:0] T7622;
  wire T4913;
  wire T4914;
  wire[3:0] T7623;
  wire T7624;
  wire[16:0] T4915;
  wire[16:0] T7625;
  wire[12:0] T4916;
  wire[3:0] T7626;
  wire T7627;
  wire T4917;
  wire T4918;
  wire[16:0] T4919;
  wire[16:0] T7628;
  wire[11:0] T4920;
  wire[11:0] T4921;
  wire[11:0] T7629;
  wire T4922;
  wire T4923;
  wire[4:0] T7630;
  wire T7631;
  wire[16:0] T4924;
  wire[16:0] T7632;
  wire[11:0] T4925;
  wire[4:0] T7633;
  wire T7634;
  wire T4926;
  wire T4927;
  wire[16:0] T4928;
  wire[16:0] T7635;
  wire[10:0] T4929;
  wire[10:0] T4930;
  wire[10:0] T7636;
  wire T4931;
  wire T4932;
  wire[5:0] T7637;
  wire T7638;
  wire[16:0] T4933;
  wire[16:0] T7639;
  wire[10:0] T4934;
  wire[5:0] T7640;
  wire T7641;
  wire T4935;
  wire T4936;
  wire[16:0] T4937;
  wire[16:0] T7642;
  wire[9:0] T4938;
  wire[9:0] T4939;
  wire[9:0] T7643;
  wire T4940;
  wire T4941;
  wire[6:0] T7644;
  wire T7645;
  wire[16:0] T4942;
  wire[16:0] T7646;
  wire[9:0] T4943;
  wire[6:0] T7647;
  wire T7648;
  wire T4944;
  wire T4945;
  wire[16:0] T4946;
  wire[16:0] T7649;
  wire[8:0] T4947;
  wire[8:0] T4948;
  wire[8:0] T7650;
  wire T4949;
  wire T4950;
  wire[7:0] T7651;
  wire T7652;
  wire[16:0] T4951;
  wire[16:0] T7653;
  wire[8:0] T4952;
  wire[7:0] T7654;
  wire T7655;
  wire T4953;
  wire T4954;
  wire[16:0] T4955;
  wire[16:0] T7656;
  wire[7:0] T4956;
  wire[7:0] T4957;
  wire[7:0] T7657;
  wire T4958;
  wire T4959;
  wire[8:0] T7658;
  wire T7659;
  wire[16:0] T4960;
  wire[16:0] T7660;
  wire[7:0] T4961;
  wire[8:0] T7661;
  wire T7662;
  wire T4962;
  wire T4963;
  wire[16:0] T4964;
  wire[16:0] T7663;
  wire[6:0] T4965;
  wire[6:0] T4966;
  wire[6:0] T7664;
  wire T4967;
  wire T4968;
  wire[9:0] T7665;
  wire T7666;
  wire[16:0] T4969;
  wire[16:0] T7667;
  wire[6:0] T4970;
  wire[9:0] T7668;
  wire T7669;
  wire T4971;
  wire T4972;
  wire[16:0] T4973;
  wire[16:0] T7670;
  wire[5:0] T4974;
  wire[5:0] T4975;
  wire[5:0] T7671;
  wire T4976;
  wire T4977;
  wire[10:0] T7672;
  wire T7673;
  wire[16:0] T4978;
  wire[16:0] T7674;
  wire[5:0] T4979;
  wire[10:0] T7675;
  wire T7676;
  wire T4980;
  wire T4981;
  wire[16:0] T4982;
  wire[16:0] T7677;
  wire[4:0] T4983;
  wire[4:0] T4984;
  wire[4:0] T7678;
  wire T4985;
  wire T4986;
  wire[11:0] T7679;
  wire T7680;
  wire[16:0] T4987;
  wire[16:0] T7681;
  wire[4:0] T4988;
  wire[11:0] T7682;
  wire T7683;
  wire T4989;
  wire T4990;
  wire[16:0] T4991;
  wire[16:0] T7684;
  wire[3:0] T4992;
  wire[3:0] T4993;
  wire[3:0] T7685;
  wire T4994;
  wire T4995;
  wire[12:0] T7686;
  wire T7687;
  wire[16:0] T4996;
  wire[16:0] T7688;
  wire[3:0] T4997;
  wire[12:0] T7689;
  wire T7690;
  wire T4998;
  wire T4999;
  wire[16:0] T5000;
  wire[16:0] T7691;
  wire[2:0] T5001;
  wire[2:0] T5002;
  wire[2:0] T7692;
  wire T5003;
  wire T5004;
  wire[13:0] T7693;
  wire T7694;
  wire[16:0] T5005;
  wire[16:0] T7695;
  wire[2:0] T5006;
  wire[13:0] T7696;
  wire T7697;
  wire T5007;
  wire T5008;
  wire[16:0] T5009;
  wire[16:0] T7698;
  wire[1:0] T5010;
  wire[1:0] T5011;
  wire[1:0] T7699;
  wire T5012;
  wire T5013;
  wire[14:0] T7700;
  wire T7701;
  wire[16:0] T5014;
  wire[16:0] T7702;
  wire[1:0] T5015;
  wire[14:0] T7703;
  wire T7704;
  wire T5016;
  wire T5017;
  wire[63:0] ConfigurationModule_io_out;
  wire[63:0] ConfigurationModule_1_io_out;
  wire[63:0] ConfigurationModule_2_io_out;
  wire[63:0] ConfigurationModule_3_io_out;
  wire[63:0] ConfigurationModule_4_io_out;
  wire[63:0] ConfigurationModule_5_io_out;
  wire[63:0] ConfigurationModule_6_io_out;
  wire[63:0] ConfigurationModule_7_io_out;
  wire[63:0] ConfigurationModule_8_io_out;
  wire[63:0] ConfigurationModule_9_io_out;
  wire[63:0] ConfigurationModule_10_io_out;
  wire[63:0] ConfigurationModule_11_io_out;
  wire[63:0] ConfigurationModule_12_io_out;
  wire[63:0] ConfigurationModule_13_io_out;
  wire[63:0] ConfigurationModule_14_io_out;
  wire[63:0] ConfigurationModule_15_io_out;
  wire[63:0] ConfigurationModule_16_io_out;
  wire[63:0] ConfigurationModule_17_io_out;
  wire[63:0] ConfigurationModule_18_io_out;
  wire[63:0] ConfigurationModule_19_io_out;
  wire[63:0] ConfigurationModule_20_io_out;
  wire[63:0] ConfigurationModule_21_io_out;
  wire[63:0] ConfigurationModule_22_io_out;
  wire[63:0] ConfigurationModule_23_io_out;
  wire[1:0] GWireModule_io_G_out;
  wire[1:0] GWireModule_1_io_G_out;
  wire[1:0] GWireModule_2_io_G_out;
  wire[1:0] GWireModule_3_io_G_out;
  wire[1:0] LoopWireBlackBox_out;
  wire[1:0] LoopWireBlackBox_1_out;
  wire[1:0] LoopWireBlackBox_2_out;
  wire[1:0] LoopWireBlackBox_3_out;
  wire[1:0] LoopWireBlackBox_4_out;
  wire[1:0] LoopWireBlackBox_5_out;
  wire[1:0] LoopWireBlackBox_6_out;
  wire[1:0] LoopWireBlackBox_7_out;
  wire[1:0] LoopWireBlackBox_8_out;
  wire[1:0] LoopWireBlackBox_9_out;
  wire[1:0] LoopWireBlackBox_10_out;
  wire[1:0] LoopWireBlackBox_11_out;
  wire[1:0] LoopWireBlackBox_12_out;
  wire[1:0] LoopWireBlackBox_13_out;
  wire[1:0] LoopWireBlackBox_14_out;
  wire[1:0] LoopWireBlackBox_15_out;
  wire[1:0] LoopWireBlackBox_16_out;
  wire[1:0] LoopWireBlackBox_17_out;
  wire[1:0] LoopWireBlackBox_18_out;
  wire[1:0] LoopWireBlackBox_19_out;
  wire[1:0] LoopWireBlackBox_20_out;
  wire[1:0] LoopWireBlackBox_21_out;
  wire[1:0] LoopWireBlackBox_22_out;
  wire[1:0] LoopWireBlackBox_23_out;
  wire[1:0] LoopWireBlackBox_24_out;
  wire[1:0] LoopWireBlackBox_25_out;
  wire[1:0] LoopWireBlackBox_26_out;
  wire[1:0] LoopWireBlackBox_27_out;
  wire[1:0] LoopWireBlackBox_28_out;
  wire[1:0] LoopWireBlackBox_29_out;
  wire[1:0] LoopWireBlackBox_30_out;
  wire[1:0] LoopWireBlackBox_31_out;
  wire[1:0] LoopWireBlackBox_32_out;
  wire[1:0] LoopWireBlackBox_33_out;
  wire[1:0] LoopWireBlackBox_34_out;
  wire[1:0] LoopWireBlackBox_35_out;
  wire[1:0] LoopWireBlackBox_36_out;
  wire[1:0] ControlBlockModule_io_Hdir;
  wire ControlBlockModule_io_store_transfer_access;
  wire ControlBlockModule_io_mem_D_or_Z;
  wire LogicBlockModule_io_shift_X_out_2;
  wire LogicBlockModule_io_shift_X_out_1;
  wire LogicBlockModule_io_shift_X_out_0;
  wire LogicBlockModule_io_shift_carry_out;
  wire LogicBlockModule_io_carry_out;
  wire[1:0] LogicBlockModule_io_mem_bus_out;
  wire[1:0] LogicBlockModule_io_V_wire_out;
  wire[1:0] LogicBlockModule_io_H_wire_out;
  wire[1:0] LogicBlockModule_io_G_wire_out;
  wire[2:0] LogicBlockModule_io_config_G_out;
  wire[4:0] LogicBlockModule_io_config_V_out;
  wire LogicBlockModule_1_io_shift_X_out_2;
  wire LogicBlockModule_1_io_shift_X_out_1;
  wire LogicBlockModule_1_io_shift_X_out_0;
  wire LogicBlockModule_1_io_shift_carry_out;
  wire LogicBlockModule_1_io_carry_out;
  wire[1:0] LogicBlockModule_1_io_mem_bus_out;
  wire[1:0] LogicBlockModule_1_io_V_wire_out;
  wire[1:0] LogicBlockModule_1_io_H_wire_out;
  wire[1:0] LogicBlockModule_1_io_G_wire_out;
  wire[2:0] LogicBlockModule_1_io_config_G_out;
  wire[4:0] LogicBlockModule_1_io_config_V_out;
  wire LogicBlockModule_2_io_shift_X_out_2;
  wire LogicBlockModule_2_io_shift_X_out_1;
  wire LogicBlockModule_2_io_shift_X_out_0;
  wire LogicBlockModule_2_io_shift_carry_out;
  wire LogicBlockModule_2_io_carry_out;
  wire[1:0] LogicBlockModule_2_io_mem_bus_out;
  wire[1:0] LogicBlockModule_2_io_V_wire_out;
  wire[1:0] LogicBlockModule_2_io_H_wire_out;
  wire[1:0] LogicBlockModule_2_io_G_wire_out;
  wire[2:0] LogicBlockModule_2_io_config_G_out;
  wire[4:0] LogicBlockModule_2_io_config_V_out;
  wire LogicBlockModule_3_io_shift_X_out_2;
  wire LogicBlockModule_3_io_shift_X_out_1;
  wire LogicBlockModule_3_io_shift_X_out_0;
  wire LogicBlockModule_3_io_shift_carry_out;
  wire LogicBlockModule_3_io_carry_out;
  wire[1:0] LogicBlockModule_3_io_mem_bus_out;
  wire[1:0] LogicBlockModule_3_io_V_wire_out;
  wire[1:0] LogicBlockModule_3_io_H_wire_out;
  wire[1:0] LogicBlockModule_3_io_G_wire_out;
  wire[2:0] LogicBlockModule_3_io_config_G_out;
  wire[4:0] LogicBlockModule_3_io_config_V_out;
  wire LogicBlockModule_4_io_shift_X_out_2;
  wire LogicBlockModule_4_io_shift_X_out_1;
  wire LogicBlockModule_4_io_shift_X_out_0;
  wire LogicBlockModule_4_io_shift_carry_out;
  wire LogicBlockModule_4_io_carry_out;
  wire[1:0] LogicBlockModule_4_io_mem_bus_out;
  wire[1:0] LogicBlockModule_4_io_V_wire_out;
  wire[1:0] LogicBlockModule_4_io_H_wire_out;
  wire[1:0] LogicBlockModule_4_io_G_wire_out;
  wire[2:0] LogicBlockModule_4_io_config_G_out;
  wire[4:0] LogicBlockModule_4_io_config_V_out;
  wire LogicBlockModule_5_io_shift_X_out_2;
  wire LogicBlockModule_5_io_shift_X_out_1;
  wire LogicBlockModule_5_io_shift_X_out_0;
  wire LogicBlockModule_5_io_shift_carry_out;
  wire LogicBlockModule_5_io_carry_out;
  wire[1:0] LogicBlockModule_5_io_mem_bus_out;
  wire[1:0] LogicBlockModule_5_io_V_wire_out;
  wire[1:0] LogicBlockModule_5_io_H_wire_out;
  wire[1:0] LogicBlockModule_5_io_G_wire_out;
  wire[2:0] LogicBlockModule_5_io_config_G_out;
  wire[4:0] LogicBlockModule_5_io_config_V_out;
  wire LogicBlockModule_6_io_shift_X_out_2;
  wire LogicBlockModule_6_io_shift_X_out_1;
  wire LogicBlockModule_6_io_shift_X_out_0;
  wire LogicBlockModule_6_io_shift_carry_out;
  wire LogicBlockModule_6_io_carry_out;
  wire[1:0] LogicBlockModule_6_io_mem_bus_out;
  wire[1:0] LogicBlockModule_6_io_V_wire_out;
  wire[1:0] LogicBlockModule_6_io_H_wire_out;
  wire[1:0] LogicBlockModule_6_io_G_wire_out;
  wire[2:0] LogicBlockModule_6_io_config_G_out;
  wire[4:0] LogicBlockModule_6_io_config_V_out;
  wire LogicBlockModule_7_io_shift_X_out_2;
  wire LogicBlockModule_7_io_shift_X_out_1;
  wire LogicBlockModule_7_io_shift_X_out_0;
  wire LogicBlockModule_7_io_shift_carry_out;
  wire LogicBlockModule_7_io_carry_out;
  wire[1:0] LogicBlockModule_7_io_mem_bus_out;
  wire[1:0] LogicBlockModule_7_io_V_wire_out;
  wire[1:0] LogicBlockModule_7_io_H_wire_out;
  wire[1:0] LogicBlockModule_7_io_G_wire_out;
  wire[2:0] LogicBlockModule_7_io_config_G_out;
  wire[4:0] LogicBlockModule_7_io_config_V_out;
  wire LogicBlockModule_8_io_shift_X_out_2;
  wire LogicBlockModule_8_io_shift_X_out_1;
  wire LogicBlockModule_8_io_shift_X_out_0;
  wire LogicBlockModule_8_io_shift_carry_out;
  wire LogicBlockModule_8_io_carry_out;
  wire[1:0] LogicBlockModule_8_io_mem_bus_out;
  wire[1:0] LogicBlockModule_8_io_V_wire_out;
  wire[1:0] LogicBlockModule_8_io_H_wire_out;
  wire[1:0] LogicBlockModule_8_io_G_wire_out;
  wire[2:0] LogicBlockModule_8_io_config_G_out;
  wire[4:0] LogicBlockModule_8_io_config_V_out;
  wire LogicBlockModule_9_io_shift_X_out_2;
  wire LogicBlockModule_9_io_shift_X_out_1;
  wire LogicBlockModule_9_io_shift_X_out_0;
  wire LogicBlockModule_9_io_shift_carry_out;
  wire LogicBlockModule_9_io_carry_out;
  wire[1:0] LogicBlockModule_9_io_mem_bus_out;
  wire[1:0] LogicBlockModule_9_io_V_wire_out;
  wire[1:0] LogicBlockModule_9_io_H_wire_out;
  wire[1:0] LogicBlockModule_9_io_G_wire_out;
  wire[2:0] LogicBlockModule_9_io_config_G_out;
  wire[4:0] LogicBlockModule_9_io_config_V_out;
  wire LogicBlockModule_10_io_shift_X_out_2;
  wire LogicBlockModule_10_io_shift_X_out_1;
  wire LogicBlockModule_10_io_shift_X_out_0;
  wire LogicBlockModule_10_io_shift_carry_out;
  wire LogicBlockModule_10_io_carry_out;
  wire[1:0] LogicBlockModule_10_io_mem_bus_out;
  wire[1:0] LogicBlockModule_10_io_V_wire_out;
  wire[1:0] LogicBlockModule_10_io_H_wire_out;
  wire[1:0] LogicBlockModule_10_io_G_wire_out;
  wire[2:0] LogicBlockModule_10_io_config_G_out;
  wire[4:0] LogicBlockModule_10_io_config_V_out;
  wire LogicBlockModule_11_io_shift_X_out_2;
  wire LogicBlockModule_11_io_shift_X_out_1;
  wire LogicBlockModule_11_io_shift_X_out_0;
  wire LogicBlockModule_11_io_shift_carry_out;
  wire LogicBlockModule_11_io_carry_out;
  wire[1:0] LogicBlockModule_11_io_mem_bus_out;
  wire[1:0] LogicBlockModule_11_io_V_wire_out;
  wire[1:0] LogicBlockModule_11_io_H_wire_out;
  wire[1:0] LogicBlockModule_11_io_G_wire_out;
  wire[2:0] LogicBlockModule_11_io_config_G_out;
  wire[4:0] LogicBlockModule_11_io_config_V_out;
  wire LogicBlockModule_12_io_shift_X_out_2;
  wire LogicBlockModule_12_io_shift_X_out_1;
  wire LogicBlockModule_12_io_shift_X_out_0;
  wire LogicBlockModule_12_io_shift_carry_out;
  wire LogicBlockModule_12_io_carry_out;
  wire[1:0] LogicBlockModule_12_io_mem_bus_out;
  wire[1:0] LogicBlockModule_12_io_V_wire_out;
  wire[1:0] LogicBlockModule_12_io_H_wire_out;
  wire[1:0] LogicBlockModule_12_io_G_wire_out;
  wire[2:0] LogicBlockModule_12_io_config_G_out;
  wire[4:0] LogicBlockModule_12_io_config_V_out;
  wire LogicBlockModule_13_io_shift_X_out_2;
  wire LogicBlockModule_13_io_shift_X_out_1;
  wire LogicBlockModule_13_io_shift_X_out_0;
  wire LogicBlockModule_13_io_shift_carry_out;
  wire LogicBlockModule_13_io_carry_out;
  wire[1:0] LogicBlockModule_13_io_mem_bus_out;
  wire[1:0] LogicBlockModule_13_io_V_wire_out;
  wire[1:0] LogicBlockModule_13_io_H_wire_out;
  wire[1:0] LogicBlockModule_13_io_G_wire_out;
  wire[2:0] LogicBlockModule_13_io_config_G_out;
  wire[4:0] LogicBlockModule_13_io_config_V_out;
  wire LogicBlockModule_14_io_shift_X_out_2;
  wire LogicBlockModule_14_io_shift_X_out_1;
  wire LogicBlockModule_14_io_shift_X_out_0;
  wire LogicBlockModule_14_io_shift_carry_out;
  wire LogicBlockModule_14_io_carry_out;
  wire[1:0] LogicBlockModule_14_io_mem_bus_out;
  wire[1:0] LogicBlockModule_14_io_V_wire_out;
  wire[1:0] LogicBlockModule_14_io_H_wire_out;
  wire[1:0] LogicBlockModule_14_io_G_wire_out;
  wire[2:0] LogicBlockModule_14_io_config_G_out;
  wire[4:0] LogicBlockModule_14_io_config_V_out;
  wire LogicBlockModule_15_io_shift_X_out_2;
  wire LogicBlockModule_15_io_shift_X_out_1;
  wire LogicBlockModule_15_io_shift_X_out_0;
  wire LogicBlockModule_15_io_shift_carry_out;
  wire LogicBlockModule_15_io_carry_out;
  wire[1:0] LogicBlockModule_15_io_mem_bus_out;
  wire[1:0] LogicBlockModule_15_io_V_wire_out;
  wire[1:0] LogicBlockModule_15_io_H_wire_out;
  wire[1:0] LogicBlockModule_15_io_G_wire_out;
  wire[2:0] LogicBlockModule_15_io_config_G_out;
  wire[4:0] LogicBlockModule_15_io_config_V_out;
  wire LogicBlockModule_16_io_shift_X_out_2;
  wire LogicBlockModule_16_io_shift_X_out_1;
  wire LogicBlockModule_16_io_shift_X_out_0;
  wire LogicBlockModule_16_io_shift_carry_out;
  wire LogicBlockModule_16_io_carry_out;
  wire[1:0] LogicBlockModule_16_io_mem_bus_out;
  wire[1:0] LogicBlockModule_16_io_V_wire_out;
  wire[1:0] LogicBlockModule_16_io_H_wire_out;
  wire[1:0] LogicBlockModule_16_io_G_wire_out;
  wire[2:0] LogicBlockModule_16_io_config_G_out;
  wire[4:0] LogicBlockModule_16_io_config_V_out;
  wire LogicBlockModule_17_io_shift_X_out_2;
  wire LogicBlockModule_17_io_shift_X_out_1;
  wire LogicBlockModule_17_io_shift_X_out_0;
  wire LogicBlockModule_17_io_shift_carry_out;
  wire LogicBlockModule_17_io_carry_out;
  wire[1:0] LogicBlockModule_17_io_mem_bus_out;
  wire[1:0] LogicBlockModule_17_io_V_wire_out;
  wire[1:0] LogicBlockModule_17_io_H_wire_out;
  wire[1:0] LogicBlockModule_17_io_G_wire_out;
  wire[2:0] LogicBlockModule_17_io_config_G_out;
  wire[4:0] LogicBlockModule_17_io_config_V_out;
  wire LogicBlockModule_18_io_shift_X_out_2;
  wire LogicBlockModule_18_io_shift_X_out_1;
  wire LogicBlockModule_18_io_shift_X_out_0;
  wire LogicBlockModule_18_io_shift_carry_out;
  wire LogicBlockModule_18_io_carry_out;
  wire[1:0] LogicBlockModule_18_io_mem_bus_out;
  wire[1:0] LogicBlockModule_18_io_V_wire_out;
  wire[1:0] LogicBlockModule_18_io_H_wire_out;
  wire[1:0] LogicBlockModule_18_io_G_wire_out;
  wire[2:0] LogicBlockModule_18_io_config_G_out;
  wire[4:0] LogicBlockModule_18_io_config_V_out;
  wire LogicBlockModule_19_io_shift_X_out_2;
  wire LogicBlockModule_19_io_shift_X_out_1;
  wire LogicBlockModule_19_io_shift_X_out_0;
  wire LogicBlockModule_19_io_shift_carry_out;
  wire LogicBlockModule_19_io_carry_out;
  wire[1:0] LogicBlockModule_19_io_mem_bus_out;
  wire[1:0] LogicBlockModule_19_io_V_wire_out;
  wire[1:0] LogicBlockModule_19_io_H_wire_out;
  wire[1:0] LogicBlockModule_19_io_G_wire_out;
  wire[2:0] LogicBlockModule_19_io_config_G_out;
  wire[4:0] LogicBlockModule_19_io_config_V_out;
  wire LogicBlockModule_20_io_shift_X_out_2;
  wire LogicBlockModule_20_io_shift_X_out_1;
  wire LogicBlockModule_20_io_shift_X_out_0;
  wire LogicBlockModule_20_io_shift_carry_out;
  wire LogicBlockModule_20_io_carry_out;
  wire[1:0] LogicBlockModule_20_io_mem_bus_out;
  wire[1:0] LogicBlockModule_20_io_V_wire_out;
  wire[1:0] LogicBlockModule_20_io_H_wire_out;
  wire[1:0] LogicBlockModule_20_io_G_wire_out;
  wire[2:0] LogicBlockModule_20_io_config_G_out;
  wire[4:0] LogicBlockModule_20_io_config_V_out;
  wire LogicBlockModule_21_io_shift_X_out_2;
  wire LogicBlockModule_21_io_shift_X_out_1;
  wire LogicBlockModule_21_io_shift_X_out_0;
  wire LogicBlockModule_21_io_shift_carry_out;
  wire LogicBlockModule_21_io_carry_out;
  wire[1:0] LogicBlockModule_21_io_mem_bus_out;
  wire[1:0] LogicBlockModule_21_io_V_wire_out;
  wire[1:0] LogicBlockModule_21_io_H_wire_out;
  wire[1:0] LogicBlockModule_21_io_G_wire_out;
  wire[2:0] LogicBlockModule_21_io_config_G_out;
  wire[4:0] LogicBlockModule_21_io_config_V_out;
  wire[1:0] LogicBlockModule_22_io_mem_bus_out;
  wire[1:0] LogicBlockModule_22_io_V_wire_out;
  wire[1:0] LogicBlockModule_22_io_H_wire_out;
  wire[1:0] LogicBlockModule_22_io_G_wire_out;
  wire[2:0] LogicBlockModule_22_io_config_G_out;
  wire[4:0] LogicBlockModule_22_io_config_V_out;


`ifndef SYNTHESIS
// synthesis translate_off
  assign io_mem_bus_out_23 = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = T1 ? LogicBlockModule_io_H_wire_out : 2'h0;
  assign T1 = 2'h2 == ControlBlockModule_io_Hdir;
  assign T2 = T1 ? LogicBlockModule_1_io_H_wire_out : 2'h0;
  assign T3 = T1 ? LogicBlockModule_2_io_H_wire_out : 2'h0;
  assign T4 = T1 ? LogicBlockModule_3_io_H_wire_out : 2'h0;
  assign T5 = T1 ? LogicBlockModule_4_io_H_wire_out : T6;
  assign T6 = T7 ? LogicBlockModule_io_H_wire_out : 2'h0;
  assign T7 = 2'h1 == ControlBlockModule_io_Hdir;
  assign T8 = T1 ? LogicBlockModule_5_io_H_wire_out : T9;
  assign T9 = T7 ? LogicBlockModule_1_io_H_wire_out : 2'h0;
  assign T10 = T1 ? LogicBlockModule_6_io_H_wire_out : T11;
  assign T11 = T7 ? LogicBlockModule_2_io_H_wire_out : 2'h0;
  assign T12 = T1 ? LogicBlockModule_7_io_H_wire_out : T13;
  assign T13 = T7 ? LogicBlockModule_3_io_H_wire_out : 2'h0;
  assign T14 = T1 ? LogicBlockModule_8_io_H_wire_out : T15;
  assign T15 = T7 ? LogicBlockModule_4_io_H_wire_out : T16;
  assign T16 = T17 ? LogicBlockModule_io_H_wire_out : 2'h0;
  assign T17 = 2'h0 == ControlBlockModule_io_Hdir;
  assign T18 = T1 ? LogicBlockModule_9_io_H_wire_out : T19;
  assign T19 = T7 ? LogicBlockModule_5_io_H_wire_out : T20;
  assign T20 = T17 ? LogicBlockModule_1_io_H_wire_out : 2'h0;
  assign T21 = T1 ? LogicBlockModule_10_io_H_wire_out : T22;
  assign T22 = T7 ? LogicBlockModule_6_io_H_wire_out : T23;
  assign T23 = T17 ? LogicBlockModule_2_io_H_wire_out : 2'h0;
  assign T24 = T1 ? LogicBlockModule_11_io_H_wire_out : T25;
  assign T25 = T7 ? LogicBlockModule_7_io_H_wire_out : T26;
  assign T26 = T17 ? LogicBlockModule_3_io_H_wire_out : 2'h0;
  assign T27 = T1 ? LogicBlockModule_12_io_H_wire_out : T28;
  assign T28 = T7 ? LogicBlockModule_8_io_H_wire_out : T29;
  assign T29 = T17 ? LogicBlockModule_4_io_H_wire_out : 2'h0;
  assign T30 = T1 ? LogicBlockModule_13_io_H_wire_out : T31;
  assign T31 = T7 ? LogicBlockModule_9_io_H_wire_out : T32;
  assign T32 = T17 ? LogicBlockModule_5_io_H_wire_out : 2'h0;
  assign T33 = T1 ? LogicBlockModule_14_io_H_wire_out : T34;
  assign T34 = T7 ? LogicBlockModule_10_io_H_wire_out : T35;
  assign T35 = T17 ? LogicBlockModule_6_io_H_wire_out : 2'h0;
  assign T36 = T1 ? LogicBlockModule_15_io_H_wire_out : T37;
  assign T37 = T7 ? LogicBlockModule_11_io_H_wire_out : T38;
  assign T38 = T17 ? LogicBlockModule_7_io_H_wire_out : 2'h0;
  assign T39 = T1 ? LogicBlockModule_16_io_H_wire_out : T40;
  assign T40 = T7 ? LogicBlockModule_12_io_H_wire_out : T41;
  assign T41 = T17 ? LogicBlockModule_8_io_H_wire_out : 2'h0;
  assign T42 = T1 ? LogicBlockModule_17_io_H_wire_out : T43;
  assign T43 = T7 ? LogicBlockModule_13_io_H_wire_out : T44;
  assign T44 = T17 ? LogicBlockModule_9_io_H_wire_out : 2'h0;
  assign T45 = T1 ? LogicBlockModule_18_io_H_wire_out : T46;
  assign T46 = T7 ? LogicBlockModule_14_io_H_wire_out : T47;
  assign T47 = T17 ? LogicBlockModule_10_io_H_wire_out : 2'h0;
  assign T48 = T1 ? LogicBlockModule_19_io_H_wire_out : T49;
  assign T49 = T7 ? LogicBlockModule_15_io_H_wire_out : T50;
  assign T50 = T17 ? LogicBlockModule_11_io_H_wire_out : 2'h0;
  assign T51 = T1 ? LogicBlockModule_20_io_H_wire_out : T52;
  assign T52 = T7 ? LogicBlockModule_16_io_H_wire_out : T53;
  assign T53 = T17 ? LogicBlockModule_12_io_H_wire_out : 2'h0;
  assign T54 = T1 ? LogicBlockModule_21_io_H_wire_out : T55;
  assign T55 = T7 ? LogicBlockModule_17_io_H_wire_out : T56;
  assign T56 = T17 ? LogicBlockModule_13_io_H_wire_out : 2'h0;
  assign T57 = T1 ? LogicBlockModule_22_io_H_wire_out : T58;
  assign T58 = T7 ? LogicBlockModule_18_io_H_wire_out : T59;
  assign T59 = T17 ? LogicBlockModule_14_io_H_wire_out : 2'h0;
  assign T60 = T7 ? LogicBlockModule_19_io_H_wire_out : T61;
  assign T61 = T17 ? LogicBlockModule_15_io_H_wire_out : 2'h0;
  assign T62 = T7 ? LogicBlockModule_20_io_H_wire_out : T63;
  assign T63 = T17 ? LogicBlockModule_16_io_H_wire_out : 2'h0;
  assign T64 = T7 ? LogicBlockModule_21_io_H_wire_out : T65;
  assign T65 = T17 ? LogicBlockModule_17_io_H_wire_out : 2'h0;
  assign T66 = T7 ? LogicBlockModule_22_io_H_wire_out : T67;
  assign T67 = T17 ? LogicBlockModule_18_io_H_wire_out : 2'h0;
  assign T68 = T17 ? LogicBlockModule_19_io_H_wire_out : 2'h0;
  assign T69 = T17 ? LogicBlockModule_20_io_H_wire_out : 2'h0;
  assign T70 = T17 ? LogicBlockModule_21_io_H_wire_out : 2'h0;
  assign T71 = T17 ? LogicBlockModule_22_io_H_wire_out : 2'h0;
  assign G_wire_below_en_3 = T5018;
  assign T5018 = T72[5'h16:1'h0];
  assign T72 = T366 ? T359 : T5019;
  assign T5019 = {1'h0, T73};
  assign T73 = T354 ? T347 : T5020;
  assign T5020 = {1'h0, T74};
  assign T74 = T342 ? T335 : T5021;
  assign T5021 = {1'h0, T75};
  assign T75 = T330 ? T323 : T5022;
  assign T5022 = {1'h0, T76};
  assign T76 = T318 ? T311 : T5023;
  assign T5023 = {1'h0, T77};
  assign T77 = T306 ? T299 : T5024;
  assign T5024 = {1'h0, T78};
  assign T78 = T294 ? T287 : T5025;
  assign T5025 = {1'h0, T79};
  assign T79 = T282 ? T275 : T5026;
  assign T5026 = {1'h0, T80};
  assign T80 = T270 ? T263 : T5027;
  assign T5027 = {1'h0, T81};
  assign T81 = T258 ? T251 : T5028;
  assign T5028 = {1'h0, T82};
  assign T82 = T246 ? T239 : T5029;
  assign T5029 = {1'h0, T83};
  assign T83 = T234 ? T227 : T5030;
  assign T5030 = {1'h0, T84};
  assign T84 = T222 ? T215 : T5031;
  assign T5031 = {1'h0, T85};
  assign T85 = T210 ? T203 : T5032;
  assign T5032 = {1'h0, T86};
  assign T86 = T198 ? T191 : T5033;
  assign T5033 = {1'h0, T87};
  assign T87 = T186 ? T179 : T5034;
  assign T5034 = {1'h0, T88};
  assign T88 = T174 ? T167 : T5035;
  assign T5035 = {1'h0, T89};
  assign T89 = T162 ? T155 : T5036;
  assign T5036 = {1'h0, T90};
  assign T90 = T150 ? T143 : T5037;
  assign T5037 = {1'h0, T91};
  assign T91 = T138 ? T131 : T5038;
  assign T5038 = {1'h0, T92};
  assign T92 = T126 ? T119 : T5039;
  assign T5039 = {1'h0, T93};
  assign T93 = T114 ? T107 : T5040;
  assign T5040 = {1'h0, T94};
  assign T94 = T102 ? T95 : 2'h0;
  assign T95 = T100 | T96;
  assign T96 = T5041 & T97;
  assign T97 = 2'h1;
  assign T5041 = T98 ? 2'h3 : 2'h0;
  assign T98 = T99;
  assign T99 = 1'h1;
  assign T100 = 2'h0 & T101;
  assign T101 = ~ T97;
  assign T102 = T105 & T103;
  assign T103 = 2'h0 == T104;
  assign T104 = LogicBlockModule_io_config_G_out[1'h1:1'h0];
  assign T105 = T106;
  assign T106 = LogicBlockModule_io_config_G_out[2'h2];
  assign T107 = T112 | T108;
  assign T108 = T5042 & T109;
  assign T109 = 3'h2;
  assign T5042 = T110 ? 3'h7 : 3'h0;
  assign T110 = T111;
  assign T111 = 1'h1;
  assign T112 = T5043 & T113;
  assign T113 = ~ T109;
  assign T5043 = {1'h0, T94};
  assign T114 = T117 & T115;
  assign T115 = 2'h0 == T116;
  assign T116 = LogicBlockModule_1_io_config_G_out[1'h1:1'h0];
  assign T117 = T118;
  assign T118 = LogicBlockModule_1_io_config_G_out[2'h2];
  assign T119 = T124 | T120;
  assign T120 = T5044 & T121;
  assign T121 = 4'h4;
  assign T5044 = T122 ? 4'hf : 4'h0;
  assign T122 = T123;
  assign T123 = 1'h1;
  assign T124 = T5045 & T125;
  assign T125 = ~ T121;
  assign T5045 = {1'h0, T93};
  assign T126 = T129 & T127;
  assign T127 = 2'h0 == T128;
  assign T128 = LogicBlockModule_2_io_config_G_out[1'h1:1'h0];
  assign T129 = T130;
  assign T130 = LogicBlockModule_2_io_config_G_out[2'h2];
  assign T131 = T136 | T132;
  assign T132 = T5046 & T133;
  assign T133 = 5'h8;
  assign T5046 = T134 ? 5'h1f : 5'h0;
  assign T134 = T135;
  assign T135 = 1'h1;
  assign T136 = T5047 & T137;
  assign T137 = ~ T133;
  assign T5047 = {1'h0, T92};
  assign T138 = T141 & T139;
  assign T139 = 2'h0 == T140;
  assign T140 = LogicBlockModule_3_io_config_G_out[1'h1:1'h0];
  assign T141 = T142;
  assign T142 = LogicBlockModule_3_io_config_G_out[2'h2];
  assign T143 = T148 | T144;
  assign T144 = T5048 & T145;
  assign T145 = 6'h10;
  assign T5048 = T146 ? 6'h3f : 6'h0;
  assign T146 = T147;
  assign T147 = 1'h1;
  assign T148 = T5049 & T149;
  assign T149 = ~ T145;
  assign T5049 = {1'h0, T91};
  assign T150 = T153 & T151;
  assign T151 = 2'h0 == T152;
  assign T152 = LogicBlockModule_4_io_config_G_out[1'h1:1'h0];
  assign T153 = T154;
  assign T154 = LogicBlockModule_4_io_config_G_out[2'h2];
  assign T155 = T160 | T156;
  assign T156 = T5050 & T157;
  assign T157 = 7'h20;
  assign T5050 = T158 ? 7'h7f : 7'h0;
  assign T158 = T159;
  assign T159 = 1'h1;
  assign T160 = T5051 & T161;
  assign T161 = ~ T157;
  assign T5051 = {1'h0, T90};
  assign T162 = T165 & T163;
  assign T163 = 2'h0 == T164;
  assign T164 = LogicBlockModule_5_io_config_G_out[1'h1:1'h0];
  assign T165 = T166;
  assign T166 = LogicBlockModule_5_io_config_G_out[2'h2];
  assign T167 = T172 | T168;
  assign T168 = T5052 & T169;
  assign T169 = 8'h40;
  assign T5052 = T170 ? 8'hff : 8'h0;
  assign T170 = T171;
  assign T171 = 1'h1;
  assign T172 = T5053 & T173;
  assign T173 = ~ T169;
  assign T5053 = {1'h0, T89};
  assign T174 = T177 & T175;
  assign T175 = 2'h0 == T176;
  assign T176 = LogicBlockModule_6_io_config_G_out[1'h1:1'h0];
  assign T177 = T178;
  assign T178 = LogicBlockModule_6_io_config_G_out[2'h2];
  assign T179 = T184 | T180;
  assign T180 = T5054 & T181;
  assign T181 = 9'h80;
  assign T5054 = T182 ? 9'h1ff : 9'h0;
  assign T182 = T183;
  assign T183 = 1'h1;
  assign T184 = T5055 & T185;
  assign T185 = ~ T181;
  assign T5055 = {1'h0, T88};
  assign T186 = T189 & T187;
  assign T187 = 2'h0 == T188;
  assign T188 = LogicBlockModule_7_io_config_G_out[1'h1:1'h0];
  assign T189 = T190;
  assign T190 = LogicBlockModule_7_io_config_G_out[2'h2];
  assign T191 = T196 | T192;
  assign T192 = T5056 & T193;
  assign T193 = 10'h100;
  assign T5056 = T194 ? 10'h3ff : 10'h0;
  assign T194 = T195;
  assign T195 = 1'h1;
  assign T196 = T5057 & T197;
  assign T197 = ~ T193;
  assign T5057 = {1'h0, T87};
  assign T198 = T201 & T199;
  assign T199 = 2'h0 == T200;
  assign T200 = LogicBlockModule_8_io_config_G_out[1'h1:1'h0];
  assign T201 = T202;
  assign T202 = LogicBlockModule_8_io_config_G_out[2'h2];
  assign T203 = T208 | T204;
  assign T204 = T5058 & T205;
  assign T205 = 11'h200;
  assign T5058 = T206 ? 11'h7ff : 11'h0;
  assign T206 = T207;
  assign T207 = 1'h1;
  assign T208 = T5059 & T209;
  assign T209 = ~ T205;
  assign T5059 = {1'h0, T86};
  assign T210 = T213 & T211;
  assign T211 = 2'h0 == T212;
  assign T212 = LogicBlockModule_9_io_config_G_out[1'h1:1'h0];
  assign T213 = T214;
  assign T214 = LogicBlockModule_9_io_config_G_out[2'h2];
  assign T215 = T220 | T216;
  assign T216 = T5060 & T217;
  assign T217 = 12'h400;
  assign T5060 = T218 ? 12'hfff : 12'h0;
  assign T218 = T219;
  assign T219 = 1'h1;
  assign T220 = T5061 & T221;
  assign T221 = ~ T217;
  assign T5061 = {1'h0, T85};
  assign T222 = T225 & T223;
  assign T223 = 2'h0 == T224;
  assign T224 = LogicBlockModule_10_io_config_G_out[1'h1:1'h0];
  assign T225 = T226;
  assign T226 = LogicBlockModule_10_io_config_G_out[2'h2];
  assign T227 = T232 | T228;
  assign T228 = T5062 & T229;
  assign T229 = 13'h800;
  assign T5062 = T230 ? 13'h1fff : 13'h0;
  assign T230 = T231;
  assign T231 = 1'h1;
  assign T232 = T5063 & T233;
  assign T233 = ~ T229;
  assign T5063 = {1'h0, T84};
  assign T234 = T237 & T235;
  assign T235 = 2'h0 == T236;
  assign T236 = LogicBlockModule_11_io_config_G_out[1'h1:1'h0];
  assign T237 = T238;
  assign T238 = LogicBlockModule_11_io_config_G_out[2'h2];
  assign T239 = T244 | T240;
  assign T240 = T5064 & T241;
  assign T241 = 14'h1000;
  assign T5064 = T242 ? 14'h3fff : 14'h0;
  assign T242 = T243;
  assign T243 = 1'h1;
  assign T244 = T5065 & T245;
  assign T245 = ~ T241;
  assign T5065 = {1'h0, T83};
  assign T246 = T249 & T247;
  assign T247 = 2'h0 == T248;
  assign T248 = LogicBlockModule_12_io_config_G_out[1'h1:1'h0];
  assign T249 = T250;
  assign T250 = LogicBlockModule_12_io_config_G_out[2'h2];
  assign T251 = T256 | T252;
  assign T252 = T5066 & T253;
  assign T253 = 15'h2000;
  assign T5066 = T254 ? 15'h7fff : 15'h0;
  assign T254 = T255;
  assign T255 = 1'h1;
  assign T256 = T5067 & T257;
  assign T257 = ~ T253;
  assign T5067 = {1'h0, T82};
  assign T258 = T261 & T259;
  assign T259 = 2'h0 == T260;
  assign T260 = LogicBlockModule_13_io_config_G_out[1'h1:1'h0];
  assign T261 = T262;
  assign T262 = LogicBlockModule_13_io_config_G_out[2'h2];
  assign T263 = T268 | T264;
  assign T264 = T5068 & T265;
  assign T265 = 16'h4000;
  assign T5068 = T266 ? 16'hffff : 16'h0;
  assign T266 = T267;
  assign T267 = 1'h1;
  assign T268 = T5069 & T269;
  assign T269 = ~ T265;
  assign T5069 = {1'h0, T81};
  assign T270 = T273 & T271;
  assign T271 = 2'h0 == T272;
  assign T272 = LogicBlockModule_14_io_config_G_out[1'h1:1'h0];
  assign T273 = T274;
  assign T274 = LogicBlockModule_14_io_config_G_out[2'h2];
  assign T275 = T280 | T276;
  assign T276 = T5070 & T277;
  assign T277 = 17'h8000;
  assign T5070 = T278 ? 17'h1ffff : 17'h0;
  assign T278 = T279;
  assign T279 = 1'h1;
  assign T280 = T5071 & T281;
  assign T281 = ~ T277;
  assign T5071 = {1'h0, T80};
  assign T282 = T285 & T283;
  assign T283 = 2'h0 == T284;
  assign T284 = LogicBlockModule_15_io_config_G_out[1'h1:1'h0];
  assign T285 = T286;
  assign T286 = LogicBlockModule_15_io_config_G_out[2'h2];
  assign T287 = T292 | T288;
  assign T288 = T5072 & T289;
  assign T289 = 18'h10000;
  assign T5072 = T290 ? 18'h3ffff : 18'h0;
  assign T290 = T291;
  assign T291 = 1'h1;
  assign T292 = T5073 & T293;
  assign T293 = ~ T289;
  assign T5073 = {1'h0, T79};
  assign T294 = T297 & T295;
  assign T295 = 2'h0 == T296;
  assign T296 = LogicBlockModule_16_io_config_G_out[1'h1:1'h0];
  assign T297 = T298;
  assign T298 = LogicBlockModule_16_io_config_G_out[2'h2];
  assign T299 = T304 | T300;
  assign T300 = T5074 & T301;
  assign T301 = 19'h20000;
  assign T5074 = T302 ? 19'h7ffff : 19'h0;
  assign T302 = T303;
  assign T303 = 1'h1;
  assign T304 = T5075 & T305;
  assign T305 = ~ T301;
  assign T5075 = {1'h0, T78};
  assign T306 = T309 & T307;
  assign T307 = 2'h0 == T308;
  assign T308 = LogicBlockModule_17_io_config_G_out[1'h1:1'h0];
  assign T309 = T310;
  assign T310 = LogicBlockModule_17_io_config_G_out[2'h2];
  assign T311 = T316 | T312;
  assign T312 = T5076 & T313;
  assign T313 = 20'h40000;
  assign T5076 = T314 ? 20'hfffff : 20'h0;
  assign T314 = T315;
  assign T315 = 1'h1;
  assign T316 = T5077 & T317;
  assign T317 = ~ T313;
  assign T5077 = {1'h0, T77};
  assign T318 = T321 & T319;
  assign T319 = 2'h0 == T320;
  assign T320 = LogicBlockModule_18_io_config_G_out[1'h1:1'h0];
  assign T321 = T322;
  assign T322 = LogicBlockModule_18_io_config_G_out[2'h2];
  assign T323 = T328 | T324;
  assign T324 = T5078 & T325;
  assign T325 = 21'h80000;
  assign T5078 = T326 ? 21'h1fffff : 21'h0;
  assign T326 = T327;
  assign T327 = 1'h1;
  assign T328 = T5079 & T329;
  assign T329 = ~ T325;
  assign T5079 = {1'h0, T76};
  assign T330 = T333 & T331;
  assign T331 = 2'h0 == T332;
  assign T332 = LogicBlockModule_19_io_config_G_out[1'h1:1'h0];
  assign T333 = T334;
  assign T334 = LogicBlockModule_19_io_config_G_out[2'h2];
  assign T335 = T340 | T336;
  assign T336 = T5080 & T337;
  assign T337 = 22'h100000;
  assign T5080 = T338 ? 22'h3fffff : 22'h0;
  assign T338 = T339;
  assign T339 = 1'h1;
  assign T340 = T5081 & T341;
  assign T341 = ~ T337;
  assign T5081 = {1'h0, T75};
  assign T342 = T345 & T343;
  assign T343 = 2'h0 == T344;
  assign T344 = LogicBlockModule_20_io_config_G_out[1'h1:1'h0];
  assign T345 = T346;
  assign T346 = LogicBlockModule_20_io_config_G_out[2'h2];
  assign T347 = T352 | T348;
  assign T348 = T5082 & T349;
  assign T349 = 23'h200000;
  assign T5082 = T350 ? 23'h7fffff : 23'h0;
  assign T350 = T351;
  assign T351 = 1'h1;
  assign T352 = T5083 & T353;
  assign T353 = ~ T349;
  assign T5083 = {1'h0, T74};
  assign T354 = T357 & T355;
  assign T355 = 2'h0 == T356;
  assign T356 = LogicBlockModule_21_io_config_G_out[1'h1:1'h0];
  assign T357 = T358;
  assign T358 = LogicBlockModule_21_io_config_G_out[2'h2];
  assign T359 = T364 | T360;
  assign T360 = T5084 & T361;
  assign T361 = 24'h400000;
  assign T5084 = T362 ? 24'hffffff : 24'h0;
  assign T362 = T363;
  assign T363 = 1'h1;
  assign T364 = T5085 & T365;
  assign T365 = ~ T361;
  assign T5085 = {1'h0, T73};
  assign T366 = T369 & T367;
  assign T367 = 2'h0 == T368;
  assign T368 = LogicBlockModule_22_io_config_G_out[1'h1:1'h0];
  assign T369 = T370;
  assign T370 = LogicBlockModule_22_io_config_G_out[2'h2];
  assign G_wire_outs_0 = LogicBlockModule_io_G_wire_out;
  assign G_wire_outs_1 = LogicBlockModule_1_io_G_wire_out;
  assign G_wire_outs_2 = LogicBlockModule_2_io_G_wire_out;
  assign G_wire_outs_3 = LogicBlockModule_3_io_G_wire_out;
  assign G_wire_outs_4 = LogicBlockModule_4_io_G_wire_out;
  assign G_wire_outs_5 = LogicBlockModule_5_io_G_wire_out;
  assign G_wire_outs_6 = LogicBlockModule_6_io_G_wire_out;
  assign G_wire_outs_7 = LogicBlockModule_7_io_G_wire_out;
  assign G_wire_outs_8 = LogicBlockModule_8_io_G_wire_out;
  assign G_wire_outs_9 = LogicBlockModule_9_io_G_wire_out;
  assign G_wire_outs_10 = LogicBlockModule_10_io_G_wire_out;
  assign G_wire_outs_11 = LogicBlockModule_11_io_G_wire_out;
  assign G_wire_outs_12 = LogicBlockModule_12_io_G_wire_out;
  assign G_wire_outs_13 = LogicBlockModule_13_io_G_wire_out;
  assign G_wire_outs_14 = LogicBlockModule_14_io_G_wire_out;
  assign G_wire_outs_15 = LogicBlockModule_15_io_G_wire_out;
  assign G_wire_outs_16 = LogicBlockModule_16_io_G_wire_out;
  assign G_wire_outs_17 = LogicBlockModule_17_io_G_wire_out;
  assign G_wire_outs_18 = LogicBlockModule_18_io_G_wire_out;
  assign G_wire_outs_19 = LogicBlockModule_19_io_G_wire_out;
  assign G_wire_outs_20 = LogicBlockModule_20_io_G_wire_out;
  assign G_wire_outs_21 = LogicBlockModule_21_io_G_wire_out;
  assign G_wire_outs_22 = LogicBlockModule_22_io_G_wire_out;
  assign G_wire_below_en_2 = T5086;
  assign T5086 = T371[5'h16:1'h0];
  assign T371 = T599 ? T592 : T5087;
  assign T5087 = {1'h0, T372};
  assign T372 = T590 ? T583 : T5088;
  assign T5088 = {1'h0, T373};
  assign T373 = T581 ? T574 : T5089;
  assign T5089 = {1'h0, T374};
  assign T374 = T572 ? T565 : T5090;
  assign T5090 = {1'h0, T375};
  assign T375 = T563 ? T556 : T5091;
  assign T5091 = {1'h0, T376};
  assign T376 = T554 ? T547 : T5092;
  assign T5092 = {1'h0, T377};
  assign T377 = T545 ? T538 : T5093;
  assign T5093 = {1'h0, T378};
  assign T378 = T536 ? T529 : T5094;
  assign T5094 = {1'h0, T379};
  assign T379 = T527 ? T520 : T5095;
  assign T5095 = {1'h0, T380};
  assign T380 = T518 ? T511 : T5096;
  assign T5096 = {1'h0, T381};
  assign T381 = T509 ? T502 : T5097;
  assign T5097 = {1'h0, T382};
  assign T382 = T500 ? T493 : T5098;
  assign T5098 = {1'h0, T383};
  assign T383 = T491 ? T484 : T5099;
  assign T5099 = {1'h0, T384};
  assign T384 = T482 ? T475 : T5100;
  assign T5100 = {1'h0, T385};
  assign T385 = T473 ? T466 : T5101;
  assign T5101 = {1'h0, T386};
  assign T386 = T464 ? T457 : T5102;
  assign T5102 = {1'h0, T387};
  assign T387 = T455 ? T448 : T5103;
  assign T5103 = {1'h0, T388};
  assign T388 = T446 ? T439 : T5104;
  assign T5104 = {1'h0, T389};
  assign T389 = T437 ? T430 : T5105;
  assign T5105 = {1'h0, T390};
  assign T390 = T428 ? T421 : T5106;
  assign T5106 = {1'h0, T391};
  assign T391 = T419 ? T412 : T5107;
  assign T5107 = {1'h0, T392};
  assign T392 = T410 ? T403 : T5108;
  assign T5108 = {1'h0, T393};
  assign T393 = T401 ? T394 : 2'h0;
  assign T394 = T399 | T395;
  assign T395 = T5109 & T396;
  assign T396 = 2'h1;
  assign T5109 = T397 ? 2'h3 : 2'h0;
  assign T397 = T398;
  assign T398 = 1'h1;
  assign T399 = 2'h0 & T400;
  assign T400 = ~ T396;
  assign T401 = T105 & T402;
  assign T402 = 2'h1 == T104;
  assign T403 = T408 | T404;
  assign T404 = T5110 & T405;
  assign T405 = 3'h2;
  assign T5110 = T406 ? 3'h7 : 3'h0;
  assign T406 = T407;
  assign T407 = 1'h1;
  assign T408 = T5111 & T409;
  assign T409 = ~ T405;
  assign T5111 = {1'h0, T393};
  assign T410 = T117 & T411;
  assign T411 = 2'h1 == T116;
  assign T412 = T417 | T413;
  assign T413 = T5112 & T414;
  assign T414 = 4'h4;
  assign T5112 = T415 ? 4'hf : 4'h0;
  assign T415 = T416;
  assign T416 = 1'h1;
  assign T417 = T5113 & T418;
  assign T418 = ~ T414;
  assign T5113 = {1'h0, T392};
  assign T419 = T129 & T420;
  assign T420 = 2'h1 == T128;
  assign T421 = T426 | T422;
  assign T422 = T5114 & T423;
  assign T423 = 5'h8;
  assign T5114 = T424 ? 5'h1f : 5'h0;
  assign T424 = T425;
  assign T425 = 1'h1;
  assign T426 = T5115 & T427;
  assign T427 = ~ T423;
  assign T5115 = {1'h0, T391};
  assign T428 = T141 & T429;
  assign T429 = 2'h1 == T140;
  assign T430 = T435 | T431;
  assign T431 = T5116 & T432;
  assign T432 = 6'h10;
  assign T5116 = T433 ? 6'h3f : 6'h0;
  assign T433 = T434;
  assign T434 = 1'h1;
  assign T435 = T5117 & T436;
  assign T436 = ~ T432;
  assign T5117 = {1'h0, T390};
  assign T437 = T153 & T438;
  assign T438 = 2'h1 == T152;
  assign T439 = T444 | T440;
  assign T440 = T5118 & T441;
  assign T441 = 7'h20;
  assign T5118 = T442 ? 7'h7f : 7'h0;
  assign T442 = T443;
  assign T443 = 1'h1;
  assign T444 = T5119 & T445;
  assign T445 = ~ T441;
  assign T5119 = {1'h0, T389};
  assign T446 = T165 & T447;
  assign T447 = 2'h1 == T164;
  assign T448 = T453 | T449;
  assign T449 = T5120 & T450;
  assign T450 = 8'h40;
  assign T5120 = T451 ? 8'hff : 8'h0;
  assign T451 = T452;
  assign T452 = 1'h1;
  assign T453 = T5121 & T454;
  assign T454 = ~ T450;
  assign T5121 = {1'h0, T388};
  assign T455 = T177 & T456;
  assign T456 = 2'h1 == T176;
  assign T457 = T462 | T458;
  assign T458 = T5122 & T459;
  assign T459 = 9'h80;
  assign T5122 = T460 ? 9'h1ff : 9'h0;
  assign T460 = T461;
  assign T461 = 1'h1;
  assign T462 = T5123 & T463;
  assign T463 = ~ T459;
  assign T5123 = {1'h0, T387};
  assign T464 = T189 & T465;
  assign T465 = 2'h1 == T188;
  assign T466 = T471 | T467;
  assign T467 = T5124 & T468;
  assign T468 = 10'h100;
  assign T5124 = T469 ? 10'h3ff : 10'h0;
  assign T469 = T470;
  assign T470 = 1'h1;
  assign T471 = T5125 & T472;
  assign T472 = ~ T468;
  assign T5125 = {1'h0, T386};
  assign T473 = T201 & T474;
  assign T474 = 2'h1 == T200;
  assign T475 = T480 | T476;
  assign T476 = T5126 & T477;
  assign T477 = 11'h200;
  assign T5126 = T478 ? 11'h7ff : 11'h0;
  assign T478 = T479;
  assign T479 = 1'h1;
  assign T480 = T5127 & T481;
  assign T481 = ~ T477;
  assign T5127 = {1'h0, T385};
  assign T482 = T213 & T483;
  assign T483 = 2'h1 == T212;
  assign T484 = T489 | T485;
  assign T485 = T5128 & T486;
  assign T486 = 12'h400;
  assign T5128 = T487 ? 12'hfff : 12'h0;
  assign T487 = T488;
  assign T488 = 1'h1;
  assign T489 = T5129 & T490;
  assign T490 = ~ T486;
  assign T5129 = {1'h0, T384};
  assign T491 = T225 & T492;
  assign T492 = 2'h1 == T224;
  assign T493 = T498 | T494;
  assign T494 = T5130 & T495;
  assign T495 = 13'h800;
  assign T5130 = T496 ? 13'h1fff : 13'h0;
  assign T496 = T497;
  assign T497 = 1'h1;
  assign T498 = T5131 & T499;
  assign T499 = ~ T495;
  assign T5131 = {1'h0, T383};
  assign T500 = T237 & T501;
  assign T501 = 2'h1 == T236;
  assign T502 = T507 | T503;
  assign T503 = T5132 & T504;
  assign T504 = 14'h1000;
  assign T5132 = T505 ? 14'h3fff : 14'h0;
  assign T505 = T506;
  assign T506 = 1'h1;
  assign T507 = T5133 & T508;
  assign T508 = ~ T504;
  assign T5133 = {1'h0, T382};
  assign T509 = T249 & T510;
  assign T510 = 2'h1 == T248;
  assign T511 = T516 | T512;
  assign T512 = T5134 & T513;
  assign T513 = 15'h2000;
  assign T5134 = T514 ? 15'h7fff : 15'h0;
  assign T514 = T515;
  assign T515 = 1'h1;
  assign T516 = T5135 & T517;
  assign T517 = ~ T513;
  assign T5135 = {1'h0, T381};
  assign T518 = T261 & T519;
  assign T519 = 2'h1 == T260;
  assign T520 = T525 | T521;
  assign T521 = T5136 & T522;
  assign T522 = 16'h4000;
  assign T5136 = T523 ? 16'hffff : 16'h0;
  assign T523 = T524;
  assign T524 = 1'h1;
  assign T525 = T5137 & T526;
  assign T526 = ~ T522;
  assign T5137 = {1'h0, T380};
  assign T527 = T273 & T528;
  assign T528 = 2'h1 == T272;
  assign T529 = T534 | T530;
  assign T530 = T5138 & T531;
  assign T531 = 17'h8000;
  assign T5138 = T532 ? 17'h1ffff : 17'h0;
  assign T532 = T533;
  assign T533 = 1'h1;
  assign T534 = T5139 & T535;
  assign T535 = ~ T531;
  assign T5139 = {1'h0, T379};
  assign T536 = T285 & T537;
  assign T537 = 2'h1 == T284;
  assign T538 = T543 | T539;
  assign T539 = T5140 & T540;
  assign T540 = 18'h10000;
  assign T5140 = T541 ? 18'h3ffff : 18'h0;
  assign T541 = T542;
  assign T542 = 1'h1;
  assign T543 = T5141 & T544;
  assign T544 = ~ T540;
  assign T5141 = {1'h0, T378};
  assign T545 = T297 & T546;
  assign T546 = 2'h1 == T296;
  assign T547 = T552 | T548;
  assign T548 = T5142 & T549;
  assign T549 = 19'h20000;
  assign T5142 = T550 ? 19'h7ffff : 19'h0;
  assign T550 = T551;
  assign T551 = 1'h1;
  assign T552 = T5143 & T553;
  assign T553 = ~ T549;
  assign T5143 = {1'h0, T377};
  assign T554 = T309 & T555;
  assign T555 = 2'h1 == T308;
  assign T556 = T561 | T557;
  assign T557 = T5144 & T558;
  assign T558 = 20'h40000;
  assign T5144 = T559 ? 20'hfffff : 20'h0;
  assign T559 = T560;
  assign T560 = 1'h1;
  assign T561 = T5145 & T562;
  assign T562 = ~ T558;
  assign T5145 = {1'h0, T376};
  assign T563 = T321 & T564;
  assign T564 = 2'h1 == T320;
  assign T565 = T570 | T566;
  assign T566 = T5146 & T567;
  assign T567 = 21'h80000;
  assign T5146 = T568 ? 21'h1fffff : 21'h0;
  assign T568 = T569;
  assign T569 = 1'h1;
  assign T570 = T5147 & T571;
  assign T571 = ~ T567;
  assign T5147 = {1'h0, T375};
  assign T572 = T333 & T573;
  assign T573 = 2'h1 == T332;
  assign T574 = T579 | T575;
  assign T575 = T5148 & T576;
  assign T576 = 22'h100000;
  assign T5148 = T577 ? 22'h3fffff : 22'h0;
  assign T577 = T578;
  assign T578 = 1'h1;
  assign T579 = T5149 & T580;
  assign T580 = ~ T576;
  assign T5149 = {1'h0, T374};
  assign T581 = T345 & T582;
  assign T582 = 2'h1 == T344;
  assign T583 = T588 | T584;
  assign T584 = T5150 & T585;
  assign T585 = 23'h200000;
  assign T5150 = T586 ? 23'h7fffff : 23'h0;
  assign T586 = T587;
  assign T587 = 1'h1;
  assign T588 = T5151 & T589;
  assign T589 = ~ T585;
  assign T5151 = {1'h0, T373};
  assign T590 = T357 & T591;
  assign T591 = 2'h1 == T356;
  assign T592 = T597 | T593;
  assign T593 = T5152 & T594;
  assign T594 = 24'h400000;
  assign T5152 = T595 ? 24'hffffff : 24'h0;
  assign T595 = T596;
  assign T596 = 1'h1;
  assign T597 = T5153 & T598;
  assign T598 = ~ T594;
  assign T5153 = {1'h0, T372};
  assign T599 = T369 & T600;
  assign T600 = 2'h1 == T368;
  assign G_wire_below_en_1 = T5154;
  assign T5154 = T601[5'h16:1'h0];
  assign T601 = T829 ? T822 : T5155;
  assign T5155 = {1'h0, T602};
  assign T602 = T820 ? T813 : T5156;
  assign T5156 = {1'h0, T603};
  assign T603 = T811 ? T804 : T5157;
  assign T5157 = {1'h0, T604};
  assign T604 = T802 ? T795 : T5158;
  assign T5158 = {1'h0, T605};
  assign T605 = T793 ? T786 : T5159;
  assign T5159 = {1'h0, T606};
  assign T606 = T784 ? T777 : T5160;
  assign T5160 = {1'h0, T607};
  assign T607 = T775 ? T768 : T5161;
  assign T5161 = {1'h0, T608};
  assign T608 = T766 ? T759 : T5162;
  assign T5162 = {1'h0, T609};
  assign T609 = T757 ? T750 : T5163;
  assign T5163 = {1'h0, T610};
  assign T610 = T748 ? T741 : T5164;
  assign T5164 = {1'h0, T611};
  assign T611 = T739 ? T732 : T5165;
  assign T5165 = {1'h0, T612};
  assign T612 = T730 ? T723 : T5166;
  assign T5166 = {1'h0, T613};
  assign T613 = T721 ? T714 : T5167;
  assign T5167 = {1'h0, T614};
  assign T614 = T712 ? T705 : T5168;
  assign T5168 = {1'h0, T615};
  assign T615 = T703 ? T696 : T5169;
  assign T5169 = {1'h0, T616};
  assign T616 = T694 ? T687 : T5170;
  assign T5170 = {1'h0, T617};
  assign T617 = T685 ? T678 : T5171;
  assign T5171 = {1'h0, T618};
  assign T618 = T676 ? T669 : T5172;
  assign T5172 = {1'h0, T619};
  assign T619 = T667 ? T660 : T5173;
  assign T5173 = {1'h0, T620};
  assign T620 = T658 ? T651 : T5174;
  assign T5174 = {1'h0, T621};
  assign T621 = T649 ? T642 : T5175;
  assign T5175 = {1'h0, T622};
  assign T622 = T640 ? T633 : T5176;
  assign T5176 = {1'h0, T623};
  assign T623 = T631 ? T624 : 2'h0;
  assign T624 = T629 | T625;
  assign T625 = T5177 & T626;
  assign T626 = 2'h1;
  assign T5177 = T627 ? 2'h3 : 2'h0;
  assign T627 = T628;
  assign T628 = 1'h1;
  assign T629 = 2'h0 & T630;
  assign T630 = ~ T626;
  assign T631 = T105 & T632;
  assign T632 = 2'h2 == T104;
  assign T633 = T638 | T634;
  assign T634 = T5178 & T635;
  assign T635 = 3'h2;
  assign T5178 = T636 ? 3'h7 : 3'h0;
  assign T636 = T637;
  assign T637 = 1'h1;
  assign T638 = T5179 & T639;
  assign T639 = ~ T635;
  assign T5179 = {1'h0, T623};
  assign T640 = T117 & T641;
  assign T641 = 2'h2 == T116;
  assign T642 = T647 | T643;
  assign T643 = T5180 & T644;
  assign T644 = 4'h4;
  assign T5180 = T645 ? 4'hf : 4'h0;
  assign T645 = T646;
  assign T646 = 1'h1;
  assign T647 = T5181 & T648;
  assign T648 = ~ T644;
  assign T5181 = {1'h0, T622};
  assign T649 = T129 & T650;
  assign T650 = 2'h2 == T128;
  assign T651 = T656 | T652;
  assign T652 = T5182 & T653;
  assign T653 = 5'h8;
  assign T5182 = T654 ? 5'h1f : 5'h0;
  assign T654 = T655;
  assign T655 = 1'h1;
  assign T656 = T5183 & T657;
  assign T657 = ~ T653;
  assign T5183 = {1'h0, T621};
  assign T658 = T141 & T659;
  assign T659 = 2'h2 == T140;
  assign T660 = T665 | T661;
  assign T661 = T5184 & T662;
  assign T662 = 6'h10;
  assign T5184 = T663 ? 6'h3f : 6'h0;
  assign T663 = T664;
  assign T664 = 1'h1;
  assign T665 = T5185 & T666;
  assign T666 = ~ T662;
  assign T5185 = {1'h0, T620};
  assign T667 = T153 & T668;
  assign T668 = 2'h2 == T152;
  assign T669 = T674 | T670;
  assign T670 = T5186 & T671;
  assign T671 = 7'h20;
  assign T5186 = T672 ? 7'h7f : 7'h0;
  assign T672 = T673;
  assign T673 = 1'h1;
  assign T674 = T5187 & T675;
  assign T675 = ~ T671;
  assign T5187 = {1'h0, T619};
  assign T676 = T165 & T677;
  assign T677 = 2'h2 == T164;
  assign T678 = T683 | T679;
  assign T679 = T5188 & T680;
  assign T680 = 8'h40;
  assign T5188 = T681 ? 8'hff : 8'h0;
  assign T681 = T682;
  assign T682 = 1'h1;
  assign T683 = T5189 & T684;
  assign T684 = ~ T680;
  assign T5189 = {1'h0, T618};
  assign T685 = T177 & T686;
  assign T686 = 2'h2 == T176;
  assign T687 = T692 | T688;
  assign T688 = T5190 & T689;
  assign T689 = 9'h80;
  assign T5190 = T690 ? 9'h1ff : 9'h0;
  assign T690 = T691;
  assign T691 = 1'h1;
  assign T692 = T5191 & T693;
  assign T693 = ~ T689;
  assign T5191 = {1'h0, T617};
  assign T694 = T189 & T695;
  assign T695 = 2'h2 == T188;
  assign T696 = T701 | T697;
  assign T697 = T5192 & T698;
  assign T698 = 10'h100;
  assign T5192 = T699 ? 10'h3ff : 10'h0;
  assign T699 = T700;
  assign T700 = 1'h1;
  assign T701 = T5193 & T702;
  assign T702 = ~ T698;
  assign T5193 = {1'h0, T616};
  assign T703 = T201 & T704;
  assign T704 = 2'h2 == T200;
  assign T705 = T710 | T706;
  assign T706 = T5194 & T707;
  assign T707 = 11'h200;
  assign T5194 = T708 ? 11'h7ff : 11'h0;
  assign T708 = T709;
  assign T709 = 1'h1;
  assign T710 = T5195 & T711;
  assign T711 = ~ T707;
  assign T5195 = {1'h0, T615};
  assign T712 = T213 & T713;
  assign T713 = 2'h2 == T212;
  assign T714 = T719 | T715;
  assign T715 = T5196 & T716;
  assign T716 = 12'h400;
  assign T5196 = T717 ? 12'hfff : 12'h0;
  assign T717 = T718;
  assign T718 = 1'h1;
  assign T719 = T5197 & T720;
  assign T720 = ~ T716;
  assign T5197 = {1'h0, T614};
  assign T721 = T225 & T722;
  assign T722 = 2'h2 == T224;
  assign T723 = T728 | T724;
  assign T724 = T5198 & T725;
  assign T725 = 13'h800;
  assign T5198 = T726 ? 13'h1fff : 13'h0;
  assign T726 = T727;
  assign T727 = 1'h1;
  assign T728 = T5199 & T729;
  assign T729 = ~ T725;
  assign T5199 = {1'h0, T613};
  assign T730 = T237 & T731;
  assign T731 = 2'h2 == T236;
  assign T732 = T737 | T733;
  assign T733 = T5200 & T734;
  assign T734 = 14'h1000;
  assign T5200 = T735 ? 14'h3fff : 14'h0;
  assign T735 = T736;
  assign T736 = 1'h1;
  assign T737 = T5201 & T738;
  assign T738 = ~ T734;
  assign T5201 = {1'h0, T612};
  assign T739 = T249 & T740;
  assign T740 = 2'h2 == T248;
  assign T741 = T746 | T742;
  assign T742 = T5202 & T743;
  assign T743 = 15'h2000;
  assign T5202 = T744 ? 15'h7fff : 15'h0;
  assign T744 = T745;
  assign T745 = 1'h1;
  assign T746 = T5203 & T747;
  assign T747 = ~ T743;
  assign T5203 = {1'h0, T611};
  assign T748 = T261 & T749;
  assign T749 = 2'h2 == T260;
  assign T750 = T755 | T751;
  assign T751 = T5204 & T752;
  assign T752 = 16'h4000;
  assign T5204 = T753 ? 16'hffff : 16'h0;
  assign T753 = T754;
  assign T754 = 1'h1;
  assign T755 = T5205 & T756;
  assign T756 = ~ T752;
  assign T5205 = {1'h0, T610};
  assign T757 = T273 & T758;
  assign T758 = 2'h2 == T272;
  assign T759 = T764 | T760;
  assign T760 = T5206 & T761;
  assign T761 = 17'h8000;
  assign T5206 = T762 ? 17'h1ffff : 17'h0;
  assign T762 = T763;
  assign T763 = 1'h1;
  assign T764 = T5207 & T765;
  assign T765 = ~ T761;
  assign T5207 = {1'h0, T609};
  assign T766 = T285 & T767;
  assign T767 = 2'h2 == T284;
  assign T768 = T773 | T769;
  assign T769 = T5208 & T770;
  assign T770 = 18'h10000;
  assign T5208 = T771 ? 18'h3ffff : 18'h0;
  assign T771 = T772;
  assign T772 = 1'h1;
  assign T773 = T5209 & T774;
  assign T774 = ~ T770;
  assign T5209 = {1'h0, T608};
  assign T775 = T297 & T776;
  assign T776 = 2'h2 == T296;
  assign T777 = T782 | T778;
  assign T778 = T5210 & T779;
  assign T779 = 19'h20000;
  assign T5210 = T780 ? 19'h7ffff : 19'h0;
  assign T780 = T781;
  assign T781 = 1'h1;
  assign T782 = T5211 & T783;
  assign T783 = ~ T779;
  assign T5211 = {1'h0, T607};
  assign T784 = T309 & T785;
  assign T785 = 2'h2 == T308;
  assign T786 = T791 | T787;
  assign T787 = T5212 & T788;
  assign T788 = 20'h40000;
  assign T5212 = T789 ? 20'hfffff : 20'h0;
  assign T789 = T790;
  assign T790 = 1'h1;
  assign T791 = T5213 & T792;
  assign T792 = ~ T788;
  assign T5213 = {1'h0, T606};
  assign T793 = T321 & T794;
  assign T794 = 2'h2 == T320;
  assign T795 = T800 | T796;
  assign T796 = T5214 & T797;
  assign T797 = 21'h80000;
  assign T5214 = T798 ? 21'h1fffff : 21'h0;
  assign T798 = T799;
  assign T799 = 1'h1;
  assign T800 = T5215 & T801;
  assign T801 = ~ T797;
  assign T5215 = {1'h0, T605};
  assign T802 = T333 & T803;
  assign T803 = 2'h2 == T332;
  assign T804 = T809 | T805;
  assign T805 = T5216 & T806;
  assign T806 = 22'h100000;
  assign T5216 = T807 ? 22'h3fffff : 22'h0;
  assign T807 = T808;
  assign T808 = 1'h1;
  assign T809 = T5217 & T810;
  assign T810 = ~ T806;
  assign T5217 = {1'h0, T604};
  assign T811 = T345 & T812;
  assign T812 = 2'h2 == T344;
  assign T813 = T818 | T814;
  assign T814 = T5218 & T815;
  assign T815 = 23'h200000;
  assign T5218 = T816 ? 23'h7fffff : 23'h0;
  assign T816 = T817;
  assign T817 = 1'h1;
  assign T818 = T5219 & T819;
  assign T819 = ~ T815;
  assign T5219 = {1'h0, T603};
  assign T820 = T357 & T821;
  assign T821 = 2'h2 == T356;
  assign T822 = T827 | T823;
  assign T823 = T5220 & T824;
  assign T824 = 24'h400000;
  assign T5220 = T825 ? 24'hffffff : 24'h0;
  assign T825 = T826;
  assign T826 = 1'h1;
  assign T827 = T5221 & T828;
  assign T828 = ~ T824;
  assign T5221 = {1'h0, T602};
  assign T829 = T369 & T830;
  assign T830 = 2'h2 == T368;
  assign G_wire_below_en_0 = T5222;
  assign T5222 = T831[5'h16:1'h0];
  assign T831 = T1059 ? T1052 : T5223;
  assign T5223 = {1'h0, T832};
  assign T832 = T1050 ? T1043 : T5224;
  assign T5224 = {1'h0, T833};
  assign T833 = T1041 ? T1034 : T5225;
  assign T5225 = {1'h0, T834};
  assign T834 = T1032 ? T1025 : T5226;
  assign T5226 = {1'h0, T835};
  assign T835 = T1023 ? T1016 : T5227;
  assign T5227 = {1'h0, T836};
  assign T836 = T1014 ? T1007 : T5228;
  assign T5228 = {1'h0, T837};
  assign T837 = T1005 ? T998 : T5229;
  assign T5229 = {1'h0, T838};
  assign T838 = T996 ? T989 : T5230;
  assign T5230 = {1'h0, T839};
  assign T839 = T987 ? T980 : T5231;
  assign T5231 = {1'h0, T840};
  assign T840 = T978 ? T971 : T5232;
  assign T5232 = {1'h0, T841};
  assign T841 = T969 ? T962 : T5233;
  assign T5233 = {1'h0, T842};
  assign T842 = T960 ? T953 : T5234;
  assign T5234 = {1'h0, T843};
  assign T843 = T951 ? T944 : T5235;
  assign T5235 = {1'h0, T844};
  assign T844 = T942 ? T935 : T5236;
  assign T5236 = {1'h0, T845};
  assign T845 = T933 ? T926 : T5237;
  assign T5237 = {1'h0, T846};
  assign T846 = T924 ? T917 : T5238;
  assign T5238 = {1'h0, T847};
  assign T847 = T915 ? T908 : T5239;
  assign T5239 = {1'h0, T848};
  assign T848 = T906 ? T899 : T5240;
  assign T5240 = {1'h0, T849};
  assign T849 = T897 ? T890 : T5241;
  assign T5241 = {1'h0, T850};
  assign T850 = T888 ? T881 : T5242;
  assign T5242 = {1'h0, T851};
  assign T851 = T879 ? T872 : T5243;
  assign T5243 = {1'h0, T852};
  assign T852 = T870 ? T863 : T5244;
  assign T5244 = {1'h0, T853};
  assign T853 = T861 ? T854 : 2'h0;
  assign T854 = T859 | T855;
  assign T855 = T5245 & T856;
  assign T856 = 2'h1;
  assign T5245 = T857 ? 2'h3 : 2'h0;
  assign T857 = T858;
  assign T858 = 1'h1;
  assign T859 = 2'h0 & T860;
  assign T860 = ~ T856;
  assign T861 = T105 & T862;
  assign T862 = 2'h3 == T104;
  assign T863 = T868 | T864;
  assign T864 = T5246 & T865;
  assign T865 = 3'h2;
  assign T5246 = T866 ? 3'h7 : 3'h0;
  assign T866 = T867;
  assign T867 = 1'h1;
  assign T868 = T5247 & T869;
  assign T869 = ~ T865;
  assign T5247 = {1'h0, T853};
  assign T870 = T117 & T871;
  assign T871 = 2'h3 == T116;
  assign T872 = T877 | T873;
  assign T873 = T5248 & T874;
  assign T874 = 4'h4;
  assign T5248 = T875 ? 4'hf : 4'h0;
  assign T875 = T876;
  assign T876 = 1'h1;
  assign T877 = T5249 & T878;
  assign T878 = ~ T874;
  assign T5249 = {1'h0, T852};
  assign T879 = T129 & T880;
  assign T880 = 2'h3 == T128;
  assign T881 = T886 | T882;
  assign T882 = T5250 & T883;
  assign T883 = 5'h8;
  assign T5250 = T884 ? 5'h1f : 5'h0;
  assign T884 = T885;
  assign T885 = 1'h1;
  assign T886 = T5251 & T887;
  assign T887 = ~ T883;
  assign T5251 = {1'h0, T851};
  assign T888 = T141 & T889;
  assign T889 = 2'h3 == T140;
  assign T890 = T895 | T891;
  assign T891 = T5252 & T892;
  assign T892 = 6'h10;
  assign T5252 = T893 ? 6'h3f : 6'h0;
  assign T893 = T894;
  assign T894 = 1'h1;
  assign T895 = T5253 & T896;
  assign T896 = ~ T892;
  assign T5253 = {1'h0, T850};
  assign T897 = T153 & T898;
  assign T898 = 2'h3 == T152;
  assign T899 = T904 | T900;
  assign T900 = T5254 & T901;
  assign T901 = 7'h20;
  assign T5254 = T902 ? 7'h7f : 7'h0;
  assign T902 = T903;
  assign T903 = 1'h1;
  assign T904 = T5255 & T905;
  assign T905 = ~ T901;
  assign T5255 = {1'h0, T849};
  assign T906 = T165 & T907;
  assign T907 = 2'h3 == T164;
  assign T908 = T913 | T909;
  assign T909 = T5256 & T910;
  assign T910 = 8'h40;
  assign T5256 = T911 ? 8'hff : 8'h0;
  assign T911 = T912;
  assign T912 = 1'h1;
  assign T913 = T5257 & T914;
  assign T914 = ~ T910;
  assign T5257 = {1'h0, T848};
  assign T915 = T177 & T916;
  assign T916 = 2'h3 == T176;
  assign T917 = T922 | T918;
  assign T918 = T5258 & T919;
  assign T919 = 9'h80;
  assign T5258 = T920 ? 9'h1ff : 9'h0;
  assign T920 = T921;
  assign T921 = 1'h1;
  assign T922 = T5259 & T923;
  assign T923 = ~ T919;
  assign T5259 = {1'h0, T847};
  assign T924 = T189 & T925;
  assign T925 = 2'h3 == T188;
  assign T926 = T931 | T927;
  assign T927 = T5260 & T928;
  assign T928 = 10'h100;
  assign T5260 = T929 ? 10'h3ff : 10'h0;
  assign T929 = T930;
  assign T930 = 1'h1;
  assign T931 = T5261 & T932;
  assign T932 = ~ T928;
  assign T5261 = {1'h0, T846};
  assign T933 = T201 & T934;
  assign T934 = 2'h3 == T200;
  assign T935 = T940 | T936;
  assign T936 = T5262 & T937;
  assign T937 = 11'h200;
  assign T5262 = T938 ? 11'h7ff : 11'h0;
  assign T938 = T939;
  assign T939 = 1'h1;
  assign T940 = T5263 & T941;
  assign T941 = ~ T937;
  assign T5263 = {1'h0, T845};
  assign T942 = T213 & T943;
  assign T943 = 2'h3 == T212;
  assign T944 = T949 | T945;
  assign T945 = T5264 & T946;
  assign T946 = 12'h400;
  assign T5264 = T947 ? 12'hfff : 12'h0;
  assign T947 = T948;
  assign T948 = 1'h1;
  assign T949 = T5265 & T950;
  assign T950 = ~ T946;
  assign T5265 = {1'h0, T844};
  assign T951 = T225 & T952;
  assign T952 = 2'h3 == T224;
  assign T953 = T958 | T954;
  assign T954 = T5266 & T955;
  assign T955 = 13'h800;
  assign T5266 = T956 ? 13'h1fff : 13'h0;
  assign T956 = T957;
  assign T957 = 1'h1;
  assign T958 = T5267 & T959;
  assign T959 = ~ T955;
  assign T5267 = {1'h0, T843};
  assign T960 = T237 & T961;
  assign T961 = 2'h3 == T236;
  assign T962 = T967 | T963;
  assign T963 = T5268 & T964;
  assign T964 = 14'h1000;
  assign T5268 = T965 ? 14'h3fff : 14'h0;
  assign T965 = T966;
  assign T966 = 1'h1;
  assign T967 = T5269 & T968;
  assign T968 = ~ T964;
  assign T5269 = {1'h0, T842};
  assign T969 = T249 & T970;
  assign T970 = 2'h3 == T248;
  assign T971 = T976 | T972;
  assign T972 = T5270 & T973;
  assign T973 = 15'h2000;
  assign T5270 = T974 ? 15'h7fff : 15'h0;
  assign T974 = T975;
  assign T975 = 1'h1;
  assign T976 = T5271 & T977;
  assign T977 = ~ T973;
  assign T5271 = {1'h0, T841};
  assign T978 = T261 & T979;
  assign T979 = 2'h3 == T260;
  assign T980 = T985 | T981;
  assign T981 = T5272 & T982;
  assign T982 = 16'h4000;
  assign T5272 = T983 ? 16'hffff : 16'h0;
  assign T983 = T984;
  assign T984 = 1'h1;
  assign T985 = T5273 & T986;
  assign T986 = ~ T982;
  assign T5273 = {1'h0, T840};
  assign T987 = T273 & T988;
  assign T988 = 2'h3 == T272;
  assign T989 = T994 | T990;
  assign T990 = T5274 & T991;
  assign T991 = 17'h8000;
  assign T5274 = T992 ? 17'h1ffff : 17'h0;
  assign T992 = T993;
  assign T993 = 1'h1;
  assign T994 = T5275 & T995;
  assign T995 = ~ T991;
  assign T5275 = {1'h0, T839};
  assign T996 = T285 & T997;
  assign T997 = 2'h3 == T284;
  assign T998 = T1003 | T999;
  assign T999 = T5276 & T1000;
  assign T1000 = 18'h10000;
  assign T5276 = T1001 ? 18'h3ffff : 18'h0;
  assign T1001 = T1002;
  assign T1002 = 1'h1;
  assign T1003 = T5277 & T1004;
  assign T1004 = ~ T1000;
  assign T5277 = {1'h0, T838};
  assign T1005 = T297 & T1006;
  assign T1006 = 2'h3 == T296;
  assign T1007 = T1012 | T1008;
  assign T1008 = T5278 & T1009;
  assign T1009 = 19'h20000;
  assign T5278 = T1010 ? 19'h7ffff : 19'h0;
  assign T1010 = T1011;
  assign T1011 = 1'h1;
  assign T1012 = T5279 & T1013;
  assign T1013 = ~ T1009;
  assign T5279 = {1'h0, T837};
  assign T1014 = T309 & T1015;
  assign T1015 = 2'h3 == T308;
  assign T1016 = T1021 | T1017;
  assign T1017 = T5280 & T1018;
  assign T1018 = 20'h40000;
  assign T5280 = T1019 ? 20'hfffff : 20'h0;
  assign T1019 = T1020;
  assign T1020 = 1'h1;
  assign T1021 = T5281 & T1022;
  assign T1022 = ~ T1018;
  assign T5281 = {1'h0, T836};
  assign T1023 = T321 & T1024;
  assign T1024 = 2'h3 == T320;
  assign T1025 = T1030 | T1026;
  assign T1026 = T5282 & T1027;
  assign T1027 = 21'h80000;
  assign T5282 = T1028 ? 21'h1fffff : 21'h0;
  assign T1028 = T1029;
  assign T1029 = 1'h1;
  assign T1030 = T5283 & T1031;
  assign T1031 = ~ T1027;
  assign T5283 = {1'h0, T835};
  assign T1032 = T333 & T1033;
  assign T1033 = 2'h3 == T332;
  assign T1034 = T1039 | T1035;
  assign T1035 = T5284 & T1036;
  assign T1036 = 22'h100000;
  assign T5284 = T1037 ? 22'h3fffff : 22'h0;
  assign T1037 = T1038;
  assign T1038 = 1'h1;
  assign T1039 = T5285 & T1040;
  assign T1040 = ~ T1036;
  assign T5285 = {1'h0, T834};
  assign T1041 = T345 & T1042;
  assign T1042 = 2'h3 == T344;
  assign T1043 = T1048 | T1044;
  assign T1044 = T5286 & T1045;
  assign T1045 = 23'h200000;
  assign T5286 = T1046 ? 23'h7fffff : 23'h0;
  assign T1046 = T1047;
  assign T1047 = 1'h1;
  assign T1048 = T5287 & T1049;
  assign T1049 = ~ T1045;
  assign T5287 = {1'h0, T833};
  assign T1050 = T357 & T1051;
  assign T1051 = 2'h3 == T356;
  assign T1052 = T1057 | T1053;
  assign T1053 = T5288 & T1054;
  assign T1054 = 24'h400000;
  assign T5288 = T1055 ? 24'hffffff : 24'h0;
  assign T1055 = T1056;
  assign T1056 = 1'h1;
  assign T1057 = T5289 & T1058;
  assign T1058 = ~ T1054;
  assign T5289 = {1'h0, T832};
  assign T1059 = T369 & T1060;
  assign T1060 = 2'h3 == T368;
  assign config_22 = ConfigurationModule_22_io_out;
  assign T1061 = T1062 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1062 = T1065 & T1063;
  assign T1063 = ~ T1064;
  assign T1064 = io_config_or_load;
  assign T1065 = io_row_en;
  assign T1066 = T1068 & T1067;
  assign T1067 = ~ io_config_or_load;
  assign T1068 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign G_wire_below_0 = LoopWireBlackBox_out;
  assign G_wire_below_1 = LoopWireBlackBox_1_out;
  assign G_wire_below_2 = LoopWireBlackBox_2_out;
  assign G_wire_below_3 = LoopWireBlackBox_3_out;
  assign H_wire_below_0 = LoopWireBlackBox_4_out;
  assign H_wire_below_1 = LoopWireBlackBox_5_out;
  assign H_wire_below_2 = LoopWireBlackBox_6_out;
  assign H_wire_below_3 = LoopWireBlackBox_7_out;
  assign H_wire_below_4 = LoopWireBlackBox_8_out;
  assign H_wire_below_5 = LoopWireBlackBox_9_out;
  assign H_wire_below_6 = LoopWireBlackBox_10_out;
  assign H_wire_below_7 = LoopWireBlackBox_11_out;
  assign H_wire_below_8 = LoopWireBlackBox_12_out;
  assign H_wire_below_9 = LoopWireBlackBox_13_out;
  assign H_wire_below_10 = LoopWireBlackBox_14_out;
  assign config_21 = ConfigurationModule_21_io_out;
  assign T1069 = T1070 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1070 = T1073 & T1071;
  assign T1071 = ~ T1072;
  assign T1072 = io_config_or_load;
  assign T1073 = io_row_en;
  assign T1074 = T1076 & T1075;
  assign T1075 = ~ io_config_or_load;
  assign T1076 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_11 = LoopWireBlackBox_15_out;
  assign config_20 = ConfigurationModule_20_io_out;
  assign T1077 = T1078 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1078 = T1081 & T1079;
  assign T1079 = ~ T1080;
  assign T1080 = io_config_or_load;
  assign T1081 = io_row_en;
  assign T1082 = T1084 & T1083;
  assign T1083 = ~ io_config_or_load;
  assign T1084 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_12 = LoopWireBlackBox_16_out;
  assign config_19 = ConfigurationModule_19_io_out;
  assign T1085 = T1086 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1086 = T1089 & T1087;
  assign T1087 = ~ T1088;
  assign T1088 = io_config_or_load;
  assign T1089 = io_row_en;
  assign T1090 = T1092 & T1091;
  assign T1091 = ~ io_config_or_load;
  assign T1092 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_13 = LoopWireBlackBox_17_out;
  assign config_18 = ConfigurationModule_18_io_out;
  assign T1093 = T1094 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1094 = T1097 & T1095;
  assign T1095 = ~ T1096;
  assign T1096 = io_config_or_load;
  assign T1097 = io_row_en;
  assign T1098 = T1100 & T1099;
  assign T1099 = ~ io_config_or_load;
  assign T1100 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_14 = LoopWireBlackBox_18_out;
  assign config_17 = ConfigurationModule_17_io_out;
  assign T1101 = T1102 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1102 = T1105 & T1103;
  assign T1103 = ~ T1104;
  assign T1104 = io_config_or_load;
  assign T1105 = io_row_en;
  assign T1106 = T1108 & T1107;
  assign T1107 = ~ io_config_or_load;
  assign T1108 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_15 = LoopWireBlackBox_19_out;
  assign config_16 = ConfigurationModule_16_io_out;
  assign T1109 = T1110 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1110 = T1113 & T1111;
  assign T1111 = ~ T1112;
  assign T1112 = io_config_or_load;
  assign T1113 = io_row_en;
  assign T1114 = T1116 & T1115;
  assign T1115 = ~ io_config_or_load;
  assign T1116 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_16 = LoopWireBlackBox_20_out;
  assign config_15 = ConfigurationModule_15_io_out;
  assign T1117 = T1118 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1118 = T1121 & T1119;
  assign T1119 = ~ T1120;
  assign T1120 = io_config_or_load;
  assign T1121 = io_row_en;
  assign T1122 = T1124 & T1123;
  assign T1123 = ~ io_config_or_load;
  assign T1124 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_17 = LoopWireBlackBox_21_out;
  assign config_14 = ConfigurationModule_14_io_out;
  assign T1125 = T1126 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1126 = T1129 & T1127;
  assign T1127 = ~ T1128;
  assign T1128 = io_config_or_load;
  assign T1129 = io_row_en;
  assign T1130 = T1132 & T1131;
  assign T1131 = ~ io_config_or_load;
  assign T1132 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_18 = LoopWireBlackBox_22_out;
  assign config_13 = ConfigurationModule_13_io_out;
  assign T1133 = T1134 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1134 = T1137 & T1135;
  assign T1135 = ~ T1136;
  assign T1136 = io_config_or_load;
  assign T1137 = io_row_en;
  assign T1138 = T1140 & T1139;
  assign T1139 = ~ io_config_or_load;
  assign T1140 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_19 = LoopWireBlackBox_23_out;
  assign config_12 = ConfigurationModule_12_io_out;
  assign T1141 = T1142 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1142 = T1145 & T1143;
  assign T1143 = ~ T1144;
  assign T1144 = io_config_or_load;
  assign T1145 = io_row_en;
  assign T1146 = T1148 & T1147;
  assign T1147 = ~ io_config_or_load;
  assign T1148 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_20 = LoopWireBlackBox_24_out;
  assign config_11 = ConfigurationModule_11_io_out;
  assign T1149 = T1150 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1150 = T1153 & T1151;
  assign T1151 = ~ T1152;
  assign T1152 = io_config_or_load;
  assign T1153 = io_row_en;
  assign T1154 = T1156 & T1155;
  assign T1155 = ~ io_config_or_load;
  assign T1156 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_21 = LoopWireBlackBox_25_out;
  assign config_10 = ConfigurationModule_10_io_out;
  assign T1157 = T1158 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1158 = T1161 & T1159;
  assign T1159 = ~ T1160;
  assign T1160 = io_config_or_load;
  assign T1161 = io_row_en;
  assign T1162 = T1164 & T1163;
  assign T1163 = ~ io_config_or_load;
  assign T1164 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_22 = LoopWireBlackBox_26_out;
  assign config_9 = ConfigurationModule_9_io_out;
  assign T1165 = T1166 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1166 = T1169 & T1167;
  assign T1167 = ~ T1168;
  assign T1168 = io_config_or_load;
  assign T1169 = io_row_en;
  assign T1170 = T1172 & T1171;
  assign T1171 = ~ io_config_or_load;
  assign T1172 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_23 = LoopWireBlackBox_27_out;
  assign config_8 = ConfigurationModule_8_io_out;
  assign T1173 = T1174 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1174 = T1177 & T1175;
  assign T1175 = ~ T1176;
  assign T1176 = io_config_or_load;
  assign T1177 = io_row_en;
  assign T1178 = T1180 & T1179;
  assign T1179 = ~ io_config_or_load;
  assign T1180 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_24 = LoopWireBlackBox_28_out;
  assign config_7 = ConfigurationModule_7_io_out;
  assign T1181 = T1182 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1182 = T1185 & T1183;
  assign T1183 = ~ T1184;
  assign T1184 = io_config_or_load;
  assign T1185 = io_row_en;
  assign T1186 = T1188 & T1187;
  assign T1187 = ~ io_config_or_load;
  assign T1188 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_25 = LoopWireBlackBox_29_out;
  assign config_6 = ConfigurationModule_6_io_out;
  assign T1189 = T1190 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1190 = T1193 & T1191;
  assign T1191 = ~ T1192;
  assign T1192 = io_config_or_load;
  assign T1193 = io_row_en;
  assign T1194 = T1196 & T1195;
  assign T1195 = ~ io_config_or_load;
  assign T1196 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_26 = LoopWireBlackBox_30_out;
  assign config_5 = ConfigurationModule_5_io_out;
  assign T1197 = T1198 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1198 = T1201 & T1199;
  assign T1199 = ~ T1200;
  assign T1200 = io_config_or_load;
  assign T1201 = io_row_en;
  assign T1202 = T1204 & T1203;
  assign T1203 = ~ io_config_or_load;
  assign T1204 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_27 = LoopWireBlackBox_31_out;
  assign config_4 = ConfigurationModule_4_io_out;
  assign T1205 = T1206 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1206 = T1209 & T1207;
  assign T1207 = ~ T1208;
  assign T1208 = io_config_or_load;
  assign T1209 = io_row_en;
  assign T1210 = T1212 & T1211;
  assign T1211 = ~ io_config_or_load;
  assign T1212 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_28 = LoopWireBlackBox_32_out;
  assign config_3 = ConfigurationModule_3_io_out;
  assign T1213 = T1214 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1214 = T1217 & T1215;
  assign T1215 = ~ T1216;
  assign T1216 = io_config_or_load;
  assign T1217 = io_row_en;
  assign T1218 = T1220 & T1219;
  assign T1219 = ~ io_config_or_load;
  assign T1220 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_29 = LoopWireBlackBox_33_out;
  assign config_2 = ConfigurationModule_2_io_out;
  assign T1221 = T1222 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1222 = T1225 & T1223;
  assign T1223 = ~ T1224;
  assign T1224 = io_config_or_load;
  assign T1225 = io_row_en;
  assign T1226 = T1228 & T1227;
  assign T1227 = ~ io_config_or_load;
  assign T1228 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_30 = LoopWireBlackBox_34_out;
  assign config_1 = ConfigurationModule_1_io_out;
  assign T1229 = T1230 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1230 = T1233 & T1231;
  assign T1231 = ~ T1232;
  assign T1232 = io_config_or_load;
  assign T1233 = io_row_en;
  assign T1234 = T1236 & T1235;
  assign T1235 = ~ io_config_or_load;
  assign T1236 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_31 = LoopWireBlackBox_35_out;
  assign config_0 = ConfigurationModule_io_out;
  assign T1237 = T1238 ? io_D_or_Z : ControlBlockModule_io_mem_D_or_Z;
  assign T1238 = T1241 & T1239;
  assign T1239 = ~ T1240;
  assign T1240 = io_config_or_load;
  assign T1241 = io_row_en;
  assign T1242 = T1244 & T1243;
  assign T1243 = ~ io_config_or_load;
  assign T1244 = ControlBlockModule_io_store_transfer_access & io_row_en;
  assign H_wire_below_32 = LoopWireBlackBox_36_out;
  assign config_23 = ConfigurationModule_23_io_out;
  assign T1245 = io_row_en & io_config_or_load;
  assign T1246 = io_row_en & io_config_or_load;
  assign T1247 = io_row_en & io_config_or_load;
  assign T1248 = io_row_en & io_config_or_load;
  assign T1249 = io_row_en & io_config_or_load;
  assign T1250 = io_row_en & io_config_or_load;
  assign T1251 = io_row_en & io_config_or_load;
  assign T1252 = io_row_en & io_config_or_load;
  assign T1253 = io_row_en & io_config_or_load;
  assign T1254 = io_row_en & io_config_or_load;
  assign T1255 = io_row_en & io_config_or_load;
  assign T1256 = io_row_en & io_config_or_load;
  assign T1257 = io_row_en & io_config_or_load;
  assign T1258 = io_row_en & io_config_or_load;
  assign T1259 = io_row_en & io_config_or_load;
  assign T1260 = io_row_en & io_config_or_load;
  assign T1261 = io_row_en & io_config_or_load;
  assign T1262 = io_row_en & io_config_or_load;
  assign T1263 = io_row_en & io_config_or_load;
  assign T1264 = io_row_en & io_config_or_load;
  assign T1265 = io_row_en & io_config_or_load;
  assign T1266 = io_row_en & io_config_or_load;
  assign T1267 = io_row_en & io_config_or_load;
  assign T1268 = io_row_en & io_config_or_load;
  assign io_mem_bus_out_0 = LogicBlockModule_io_mem_bus_out;
  assign io_mem_bus_out_1 = LogicBlockModule_1_io_mem_bus_out;
  assign io_mem_bus_out_2 = LogicBlockModule_2_io_mem_bus_out;
  assign io_mem_bus_out_3 = LogicBlockModule_3_io_mem_bus_out;
  assign io_mem_bus_out_4 = LogicBlockModule_4_io_mem_bus_out;
  assign io_mem_bus_out_5 = LogicBlockModule_5_io_mem_bus_out;
  assign io_mem_bus_out_6 = LogicBlockModule_6_io_mem_bus_out;
  assign io_mem_bus_out_7 = LogicBlockModule_7_io_mem_bus_out;
  assign io_mem_bus_out_8 = LogicBlockModule_8_io_mem_bus_out;
  assign io_mem_bus_out_9 = LogicBlockModule_9_io_mem_bus_out;
  assign io_mem_bus_out_10 = LogicBlockModule_10_io_mem_bus_out;
  assign io_mem_bus_out_11 = LogicBlockModule_11_io_mem_bus_out;
  assign io_mem_bus_out_12 = LogicBlockModule_12_io_mem_bus_out;
  assign io_mem_bus_out_13 = LogicBlockModule_13_io_mem_bus_out;
  assign io_mem_bus_out_14 = LogicBlockModule_14_io_mem_bus_out;
  assign io_mem_bus_out_15 = LogicBlockModule_15_io_mem_bus_out;
  assign io_mem_bus_out_16 = LogicBlockModule_16_io_mem_bus_out;
  assign io_mem_bus_out_17 = LogicBlockModule_17_io_mem_bus_out;
  assign io_mem_bus_out_18 = LogicBlockModule_18_io_mem_bus_out;
  assign io_mem_bus_out_19 = LogicBlockModule_19_io_mem_bus_out;
  assign io_mem_bus_out_20 = LogicBlockModule_20_io_mem_bus_out;
  assign io_mem_bus_out_21 = LogicBlockModule_21_io_mem_bus_out;
  assign io_mem_bus_out_22 = LogicBlockModule_22_io_mem_bus_out;
  assign io_H_wire_below_0 = H_wire_below_0;
  assign io_H_wire_below_1 = H_wire_below_1;
  assign io_H_wire_below_2 = H_wire_below_2;
  assign io_H_wire_below_3 = H_wire_below_3;
  assign io_H_wire_below_4 = H_wire_below_4;
  assign io_H_wire_below_5 = H_wire_below_5;
  assign io_H_wire_below_6 = H_wire_below_6;
  assign io_H_wire_below_7 = H_wire_below_7;
  assign io_H_wire_below_8 = H_wire_below_8;
  assign io_H_wire_below_9 = H_wire_below_9;
  assign io_H_wire_below_10 = H_wire_below_10;
  assign io_H_wire_below_11 = H_wire_below_11;
  assign io_H_wire_below_12 = H_wire_below_12;
  assign io_H_wire_below_13 = H_wire_below_13;
  assign io_H_wire_below_14 = H_wire_below_14;
  assign io_H_wire_below_15 = H_wire_below_15;
  assign io_H_wire_below_16 = H_wire_below_16;
  assign io_H_wire_below_17 = H_wire_below_17;
  assign io_H_wire_below_18 = H_wire_below_18;
  assign io_H_wire_below_19 = H_wire_below_19;
  assign io_H_wire_below_20 = H_wire_below_20;
  assign io_H_wire_below_21 = H_wire_below_21;
  assign io_H_wire_below_22 = H_wire_below_22;
  assign io_H_wire_below_23 = H_wire_below_23;
  assign io_H_wire_below_24 = H_wire_below_24;
  assign io_H_wire_below_25 = H_wire_below_25;
  assign io_H_wire_below_26 = H_wire_below_26;
  assign io_H_wire_below_27 = H_wire_below_27;
  assign io_H_wire_below_28 = H_wire_below_28;
  assign io_H_wire_below_29 = H_wire_below_29;
  assign io_H_wire_below_30 = H_wire_below_30;
  assign io_H_wire_below_31 = H_wire_below_31;
  assign io_H_wire_below_32 = H_wire_below_32;
  assign io_G_wire_below_0 = G_wire_below_0;
  assign io_G_wire_below_1 = G_wire_below_1;
  assign io_G_wire_below_2 = G_wire_below_2;
  assign io_G_wire_below_3 = G_wire_below_3;
  assign io_H_out_0 = LogicBlockModule_io_H_wire_out;
  assign io_H_out_1 = LogicBlockModule_1_io_H_wire_out;
  assign io_H_out_2 = LogicBlockModule_2_io_H_wire_out;
  assign io_H_out_3 = LogicBlockModule_3_io_H_wire_out;
  assign io_H_out_4 = LogicBlockModule_4_io_H_wire_out;
  assign io_H_out_5 = LogicBlockModule_5_io_H_wire_out;
  assign io_H_out_6 = LogicBlockModule_6_io_H_wire_out;
  assign io_H_out_7 = LogicBlockModule_7_io_H_wire_out;
  assign io_H_out_8 = LogicBlockModule_8_io_H_wire_out;
  assign io_H_out_9 = LogicBlockModule_9_io_H_wire_out;
  assign io_H_out_10 = LogicBlockModule_10_io_H_wire_out;
  assign io_H_out_11 = LogicBlockModule_11_io_H_wire_out;
  assign io_H_out_12 = LogicBlockModule_12_io_H_wire_out;
  assign io_H_out_13 = LogicBlockModule_13_io_H_wire_out;
  assign io_H_out_14 = LogicBlockModule_14_io_H_wire_out;
  assign io_H_out_15 = LogicBlockModule_15_io_H_wire_out;
  assign io_H_out_16 = LogicBlockModule_16_io_H_wire_out;
  assign io_H_out_17 = LogicBlockModule_17_io_H_wire_out;
  assign io_H_out_18 = LogicBlockModule_18_io_H_wire_out;
  assign io_H_out_19 = LogicBlockModule_19_io_H_wire_out;
  assign io_H_out_20 = LogicBlockModule_20_io_H_wire_out;
  assign io_H_out_21 = LogicBlockModule_21_io_H_wire_out;
  assign io_H_out_22 = LogicBlockModule_22_io_H_wire_out;
  assign io_V_wire_en_0 = V_wire_en_0;
  assign V_wire_en_0 = T5290;
  assign T5290 = T1269[4'hf:1'h0];
  assign T1269 = T1430 ? T1423 : T1270;
  assign T1270 = T1421 ? T1414 : T1271;
  assign T1271 = T1412 ? T1405 : T1272;
  assign T1272 = T1403 ? T1396 : T1273;
  assign T1273 = T1394 ? T1387 : T1274;
  assign T1274 = T1385 ? T1378 : T1275;
  assign T1275 = T1376 ? T1369 : T1276;
  assign T1276 = T1367 ? T1360 : T1277;
  assign T1277 = T1358 ? T1351 : T1278;
  assign T1278 = T1349 ? T1342 : T1279;
  assign T1279 = T1340 ? T1333 : T1280;
  assign T1280 = T1331 ? T1324 : T1281;
  assign T1281 = T1322 ? T1315 : T1282;
  assign T1282 = T1313 ? T1306 : T1283;
  assign T1283 = T1304 ? T1297 : T1284;
  assign T1284 = T1292 ? T1285 : 17'h0;
  assign T1285 = T1290 | T1286;
  assign T1286 = T5291 & T1287;
  assign T1287 = 17'h8000;
  assign T5291 = T1288 ? 17'h1ffff : 17'h0;
  assign T1288 = T1289;
  assign T1289 = 1'h1;
  assign T1290 = 17'h0 & T1291;
  assign T1291 = ~ T1287;
  assign T1292 = T1295 & T1293;
  assign T1293 = 4'h0 == T1294;
  assign T1294 = LogicBlockModule_io_config_V_out[2'h3:1'h0];
  assign T1295 = T1296;
  assign T1296 = LogicBlockModule_io_config_V_out[3'h4];
  assign T1297 = T1302 | T5292;
  assign T5292 = {T5294, T1298};
  assign T1298 = T5293 & T1299;
  assign T1299 = 16'h4000;
  assign T5293 = T1300 ? 16'hffff : 16'h0;
  assign T1300 = T1301;
  assign T1301 = 1'h1;
  assign T5294 = T1298[4'hf];
  assign T1302 = T1284 & T5295;
  assign T5295 = {T5296, T1303};
  assign T1303 = ~ T1299;
  assign T5296 = T1303[4'hf];
  assign T1304 = T1295 & T1305;
  assign T1305 = 4'h1 == T1294;
  assign T1306 = T1311 | T5297;
  assign T5297 = {T5299, T1307};
  assign T1307 = T5298 & T1308;
  assign T1308 = 15'h2000;
  assign T5298 = T1309 ? 15'h7fff : 15'h0;
  assign T1309 = T1310;
  assign T1310 = 1'h1;
  assign T5299 = T5300 ? 2'h3 : 2'h0;
  assign T5300 = T1307[4'he];
  assign T1311 = T1283 & T5301;
  assign T5301 = {T5302, T1312};
  assign T1312 = ~ T1308;
  assign T5302 = T5303 ? 2'h3 : 2'h0;
  assign T5303 = T1312[4'he];
  assign T1313 = T1295 & T1314;
  assign T1314 = 4'h2 == T1294;
  assign T1315 = T1320 | T5304;
  assign T5304 = {T5306, T1316};
  assign T1316 = T5305 & T1317;
  assign T1317 = 14'h1000;
  assign T5305 = T1318 ? 14'h3fff : 14'h0;
  assign T1318 = T1319;
  assign T1319 = 1'h1;
  assign T5306 = T5307 ? 3'h7 : 3'h0;
  assign T5307 = T1316[4'hd];
  assign T1320 = T1282 & T5308;
  assign T5308 = {T5309, T1321};
  assign T1321 = ~ T1317;
  assign T5309 = T5310 ? 3'h7 : 3'h0;
  assign T5310 = T1321[4'hd];
  assign T1322 = T1295 & T1323;
  assign T1323 = 4'h3 == T1294;
  assign T1324 = T1329 | T5311;
  assign T5311 = {T5313, T1325};
  assign T1325 = T5312 & T1326;
  assign T1326 = 13'h800;
  assign T5312 = T1327 ? 13'h1fff : 13'h0;
  assign T1327 = T1328;
  assign T1328 = 1'h1;
  assign T5313 = T5314 ? 4'hf : 4'h0;
  assign T5314 = T1325[4'hc];
  assign T1329 = T1281 & T5315;
  assign T5315 = {T5316, T1330};
  assign T1330 = ~ T1326;
  assign T5316 = T5317 ? 4'hf : 4'h0;
  assign T5317 = T1330[4'hc];
  assign T1331 = T1295 & T1332;
  assign T1332 = 4'h4 == T1294;
  assign T1333 = T1338 | T5318;
  assign T5318 = {T5320, T1334};
  assign T1334 = T5319 & T1335;
  assign T1335 = 12'h400;
  assign T5319 = T1336 ? 12'hfff : 12'h0;
  assign T1336 = T1337;
  assign T1337 = 1'h1;
  assign T5320 = T5321 ? 5'h1f : 5'h0;
  assign T5321 = T1334[4'hb];
  assign T1338 = T1280 & T5322;
  assign T5322 = {T5323, T1339};
  assign T1339 = ~ T1335;
  assign T5323 = T5324 ? 5'h1f : 5'h0;
  assign T5324 = T1339[4'hb];
  assign T1340 = T1295 & T1341;
  assign T1341 = 4'h5 == T1294;
  assign T1342 = T1347 | T5325;
  assign T5325 = {T5327, T1343};
  assign T1343 = T5326 & T1344;
  assign T1344 = 11'h200;
  assign T5326 = T1345 ? 11'h7ff : 11'h0;
  assign T1345 = T1346;
  assign T1346 = 1'h1;
  assign T5327 = T5328 ? 6'h3f : 6'h0;
  assign T5328 = T1343[4'ha];
  assign T1347 = T1279 & T5329;
  assign T5329 = {T5330, T1348};
  assign T1348 = ~ T1344;
  assign T5330 = T5331 ? 6'h3f : 6'h0;
  assign T5331 = T1348[4'ha];
  assign T1349 = T1295 & T1350;
  assign T1350 = 4'h6 == T1294;
  assign T1351 = T1356 | T5332;
  assign T5332 = {T5334, T1352};
  assign T1352 = T5333 & T1353;
  assign T1353 = 10'h100;
  assign T5333 = T1354 ? 10'h3ff : 10'h0;
  assign T1354 = T1355;
  assign T1355 = 1'h1;
  assign T5334 = T5335 ? 7'h7f : 7'h0;
  assign T5335 = T1352[4'h9];
  assign T1356 = T1278 & T5336;
  assign T5336 = {T5337, T1357};
  assign T1357 = ~ T1353;
  assign T5337 = T5338 ? 7'h7f : 7'h0;
  assign T5338 = T1357[4'h9];
  assign T1358 = T1295 & T1359;
  assign T1359 = 4'h7 == T1294;
  assign T1360 = T1365 | T5339;
  assign T5339 = {T5341, T1361};
  assign T1361 = T5340 & T1362;
  assign T1362 = 9'h80;
  assign T5340 = T1363 ? 9'h1ff : 9'h0;
  assign T1363 = T1364;
  assign T1364 = 1'h1;
  assign T5341 = T5342 ? 8'hff : 8'h0;
  assign T5342 = T1361[4'h8];
  assign T1365 = T1277 & T5343;
  assign T5343 = {T5344, T1366};
  assign T1366 = ~ T1362;
  assign T5344 = T5345 ? 8'hff : 8'h0;
  assign T5345 = T1366[4'h8];
  assign T1367 = T1295 & T1368;
  assign T1368 = 4'h8 == T1294;
  assign T1369 = T1374 | T5346;
  assign T5346 = {T5348, T1370};
  assign T1370 = T5347 & T1371;
  assign T1371 = 8'h40;
  assign T5347 = T1372 ? 8'hff : 8'h0;
  assign T1372 = T1373;
  assign T1373 = 1'h1;
  assign T5348 = T5349 ? 9'h1ff : 9'h0;
  assign T5349 = T1370[3'h7];
  assign T1374 = T1276 & T5350;
  assign T5350 = {T5351, T1375};
  assign T1375 = ~ T1371;
  assign T5351 = T5352 ? 9'h1ff : 9'h0;
  assign T5352 = T1375[3'h7];
  assign T1376 = T1295 & T1377;
  assign T1377 = 4'h9 == T1294;
  assign T1378 = T1383 | T5353;
  assign T5353 = {T5355, T1379};
  assign T1379 = T5354 & T1380;
  assign T1380 = 7'h20;
  assign T5354 = T1381 ? 7'h7f : 7'h0;
  assign T1381 = T1382;
  assign T1382 = 1'h1;
  assign T5355 = T5356 ? 10'h3ff : 10'h0;
  assign T5356 = T1379[3'h6];
  assign T1383 = T1275 & T5357;
  assign T5357 = {T5358, T1384};
  assign T1384 = ~ T1380;
  assign T5358 = T5359 ? 10'h3ff : 10'h0;
  assign T5359 = T1384[3'h6];
  assign T1385 = T1295 & T1386;
  assign T1386 = 4'ha == T1294;
  assign T1387 = T1392 | T5360;
  assign T5360 = {T5362, T1388};
  assign T1388 = T5361 & T1389;
  assign T1389 = 6'h10;
  assign T5361 = T1390 ? 6'h3f : 6'h0;
  assign T1390 = T1391;
  assign T1391 = 1'h1;
  assign T5362 = T5363 ? 11'h7ff : 11'h0;
  assign T5363 = T1388[3'h5];
  assign T1392 = T1274 & T5364;
  assign T5364 = {T5365, T1393};
  assign T1393 = ~ T1389;
  assign T5365 = T5366 ? 11'h7ff : 11'h0;
  assign T5366 = T1393[3'h5];
  assign T1394 = T1295 & T1395;
  assign T1395 = 4'hb == T1294;
  assign T1396 = T1401 | T5367;
  assign T5367 = {T5369, T1397};
  assign T1397 = T5368 & T1398;
  assign T1398 = 5'h8;
  assign T5368 = T1399 ? 5'h1f : 5'h0;
  assign T1399 = T1400;
  assign T1400 = 1'h1;
  assign T5369 = T5370 ? 12'hfff : 12'h0;
  assign T5370 = T1397[3'h4];
  assign T1401 = T1273 & T5371;
  assign T5371 = {T5372, T1402};
  assign T1402 = ~ T1398;
  assign T5372 = T5373 ? 12'hfff : 12'h0;
  assign T5373 = T1402[3'h4];
  assign T1403 = T1295 & T1404;
  assign T1404 = 4'hc == T1294;
  assign T1405 = T1410 | T5374;
  assign T5374 = {T5376, T1406};
  assign T1406 = T5375 & T1407;
  assign T1407 = 4'h4;
  assign T5375 = T1408 ? 4'hf : 4'h0;
  assign T1408 = T1409;
  assign T1409 = 1'h1;
  assign T5376 = T5377 ? 13'h1fff : 13'h0;
  assign T5377 = T1406[2'h3];
  assign T1410 = T1272 & T5378;
  assign T5378 = {T5379, T1411};
  assign T1411 = ~ T1407;
  assign T5379 = T5380 ? 13'h1fff : 13'h0;
  assign T5380 = T1411[2'h3];
  assign T1412 = T1295 & T1413;
  assign T1413 = 4'hd == T1294;
  assign T1414 = T1419 | T5381;
  assign T5381 = {T5383, T1415};
  assign T1415 = T5382 & T1416;
  assign T1416 = 3'h2;
  assign T5382 = T1417 ? 3'h7 : 3'h0;
  assign T1417 = T1418;
  assign T1418 = 1'h1;
  assign T5383 = T5384 ? 14'h3fff : 14'h0;
  assign T5384 = T1415[2'h2];
  assign T1419 = T1271 & T5385;
  assign T5385 = {T5386, T1420};
  assign T1420 = ~ T1416;
  assign T5386 = T5387 ? 14'h3fff : 14'h0;
  assign T5387 = T1420[2'h2];
  assign T1421 = T1295 & T1422;
  assign T1422 = 4'he == T1294;
  assign T1423 = T1428 | T5388;
  assign T5388 = {T5390, T1424};
  assign T1424 = T5389 & T1425;
  assign T1425 = 2'h1;
  assign T5389 = T1426 ? 2'h3 : 2'h0;
  assign T1426 = T1427;
  assign T1427 = 1'h1;
  assign T5390 = T5391 ? 15'h7fff : 15'h0;
  assign T5391 = T1424[1'h1];
  assign T1428 = T1270 & T5392;
  assign T5392 = {T5393, T1429};
  assign T1429 = ~ T1425;
  assign T5393 = T5394 ? 15'h7fff : 15'h0;
  assign T5394 = T1429[1'h1];
  assign T1430 = T1295 & T1431;
  assign T1431 = 4'hf == T1294;
  assign io_V_wire_en_1 = V_wire_en_1;
  assign V_wire_en_1 = T5395;
  assign T5395 = T1432[4'hf:1'h0];
  assign T1432 = T1593 ? T1586 : T1433;
  assign T1433 = T1584 ? T1577 : T1434;
  assign T1434 = T1575 ? T1568 : T1435;
  assign T1435 = T1566 ? T1559 : T1436;
  assign T1436 = T1557 ? T1550 : T1437;
  assign T1437 = T1548 ? T1541 : T1438;
  assign T1438 = T1539 ? T1532 : T1439;
  assign T1439 = T1530 ? T1523 : T1440;
  assign T1440 = T1521 ? T1514 : T1441;
  assign T1441 = T1512 ? T1505 : T1442;
  assign T1442 = T1503 ? T1496 : T1443;
  assign T1443 = T1494 ? T1487 : T1444;
  assign T1444 = T1485 ? T1478 : T1445;
  assign T1445 = T1476 ? T1469 : T1446;
  assign T1446 = T1467 ? T1460 : T1447;
  assign T1447 = T1455 ? T1448 : 17'h0;
  assign T1448 = T1453 | T1449;
  assign T1449 = T5396 & T1450;
  assign T1450 = 17'h8000;
  assign T5396 = T1451 ? 17'h1ffff : 17'h0;
  assign T1451 = T1452;
  assign T1452 = 1'h1;
  assign T1453 = 17'h0 & T1454;
  assign T1454 = ~ T1450;
  assign T1455 = T1458 & T1456;
  assign T1456 = 4'h0 == T1457;
  assign T1457 = LogicBlockModule_1_io_config_V_out[2'h3:1'h0];
  assign T1458 = T1459;
  assign T1459 = LogicBlockModule_1_io_config_V_out[3'h4];
  assign T1460 = T1465 | T5397;
  assign T5397 = {T5399, T1461};
  assign T1461 = T5398 & T1462;
  assign T1462 = 16'h4000;
  assign T5398 = T1463 ? 16'hffff : 16'h0;
  assign T1463 = T1464;
  assign T1464 = 1'h1;
  assign T5399 = T1461[4'hf];
  assign T1465 = T1447 & T5400;
  assign T5400 = {T5401, T1466};
  assign T1466 = ~ T1462;
  assign T5401 = T1466[4'hf];
  assign T1467 = T1458 & T1468;
  assign T1468 = 4'h1 == T1457;
  assign T1469 = T1474 | T5402;
  assign T5402 = {T5404, T1470};
  assign T1470 = T5403 & T1471;
  assign T1471 = 15'h2000;
  assign T5403 = T1472 ? 15'h7fff : 15'h0;
  assign T1472 = T1473;
  assign T1473 = 1'h1;
  assign T5404 = T5405 ? 2'h3 : 2'h0;
  assign T5405 = T1470[4'he];
  assign T1474 = T1446 & T5406;
  assign T5406 = {T5407, T1475};
  assign T1475 = ~ T1471;
  assign T5407 = T5408 ? 2'h3 : 2'h0;
  assign T5408 = T1475[4'he];
  assign T1476 = T1458 & T1477;
  assign T1477 = 4'h2 == T1457;
  assign T1478 = T1483 | T5409;
  assign T5409 = {T5411, T1479};
  assign T1479 = T5410 & T1480;
  assign T1480 = 14'h1000;
  assign T5410 = T1481 ? 14'h3fff : 14'h0;
  assign T1481 = T1482;
  assign T1482 = 1'h1;
  assign T5411 = T5412 ? 3'h7 : 3'h0;
  assign T5412 = T1479[4'hd];
  assign T1483 = T1445 & T5413;
  assign T5413 = {T5414, T1484};
  assign T1484 = ~ T1480;
  assign T5414 = T5415 ? 3'h7 : 3'h0;
  assign T5415 = T1484[4'hd];
  assign T1485 = T1458 & T1486;
  assign T1486 = 4'h3 == T1457;
  assign T1487 = T1492 | T5416;
  assign T5416 = {T5418, T1488};
  assign T1488 = T5417 & T1489;
  assign T1489 = 13'h800;
  assign T5417 = T1490 ? 13'h1fff : 13'h0;
  assign T1490 = T1491;
  assign T1491 = 1'h1;
  assign T5418 = T5419 ? 4'hf : 4'h0;
  assign T5419 = T1488[4'hc];
  assign T1492 = T1444 & T5420;
  assign T5420 = {T5421, T1493};
  assign T1493 = ~ T1489;
  assign T5421 = T5422 ? 4'hf : 4'h0;
  assign T5422 = T1493[4'hc];
  assign T1494 = T1458 & T1495;
  assign T1495 = 4'h4 == T1457;
  assign T1496 = T1501 | T5423;
  assign T5423 = {T5425, T1497};
  assign T1497 = T5424 & T1498;
  assign T1498 = 12'h400;
  assign T5424 = T1499 ? 12'hfff : 12'h0;
  assign T1499 = T1500;
  assign T1500 = 1'h1;
  assign T5425 = T5426 ? 5'h1f : 5'h0;
  assign T5426 = T1497[4'hb];
  assign T1501 = T1443 & T5427;
  assign T5427 = {T5428, T1502};
  assign T1502 = ~ T1498;
  assign T5428 = T5429 ? 5'h1f : 5'h0;
  assign T5429 = T1502[4'hb];
  assign T1503 = T1458 & T1504;
  assign T1504 = 4'h5 == T1457;
  assign T1505 = T1510 | T5430;
  assign T5430 = {T5432, T1506};
  assign T1506 = T5431 & T1507;
  assign T1507 = 11'h200;
  assign T5431 = T1508 ? 11'h7ff : 11'h0;
  assign T1508 = T1509;
  assign T1509 = 1'h1;
  assign T5432 = T5433 ? 6'h3f : 6'h0;
  assign T5433 = T1506[4'ha];
  assign T1510 = T1442 & T5434;
  assign T5434 = {T5435, T1511};
  assign T1511 = ~ T1507;
  assign T5435 = T5436 ? 6'h3f : 6'h0;
  assign T5436 = T1511[4'ha];
  assign T1512 = T1458 & T1513;
  assign T1513 = 4'h6 == T1457;
  assign T1514 = T1519 | T5437;
  assign T5437 = {T5439, T1515};
  assign T1515 = T5438 & T1516;
  assign T1516 = 10'h100;
  assign T5438 = T1517 ? 10'h3ff : 10'h0;
  assign T1517 = T1518;
  assign T1518 = 1'h1;
  assign T5439 = T5440 ? 7'h7f : 7'h0;
  assign T5440 = T1515[4'h9];
  assign T1519 = T1441 & T5441;
  assign T5441 = {T5442, T1520};
  assign T1520 = ~ T1516;
  assign T5442 = T5443 ? 7'h7f : 7'h0;
  assign T5443 = T1520[4'h9];
  assign T1521 = T1458 & T1522;
  assign T1522 = 4'h7 == T1457;
  assign T1523 = T1528 | T5444;
  assign T5444 = {T5446, T1524};
  assign T1524 = T5445 & T1525;
  assign T1525 = 9'h80;
  assign T5445 = T1526 ? 9'h1ff : 9'h0;
  assign T1526 = T1527;
  assign T1527 = 1'h1;
  assign T5446 = T5447 ? 8'hff : 8'h0;
  assign T5447 = T1524[4'h8];
  assign T1528 = T1440 & T5448;
  assign T5448 = {T5449, T1529};
  assign T1529 = ~ T1525;
  assign T5449 = T5450 ? 8'hff : 8'h0;
  assign T5450 = T1529[4'h8];
  assign T1530 = T1458 & T1531;
  assign T1531 = 4'h8 == T1457;
  assign T1532 = T1537 | T5451;
  assign T5451 = {T5453, T1533};
  assign T1533 = T5452 & T1534;
  assign T1534 = 8'h40;
  assign T5452 = T1535 ? 8'hff : 8'h0;
  assign T1535 = T1536;
  assign T1536 = 1'h1;
  assign T5453 = T5454 ? 9'h1ff : 9'h0;
  assign T5454 = T1533[3'h7];
  assign T1537 = T1439 & T5455;
  assign T5455 = {T5456, T1538};
  assign T1538 = ~ T1534;
  assign T5456 = T5457 ? 9'h1ff : 9'h0;
  assign T5457 = T1538[3'h7];
  assign T1539 = T1458 & T1540;
  assign T1540 = 4'h9 == T1457;
  assign T1541 = T1546 | T5458;
  assign T5458 = {T5460, T1542};
  assign T1542 = T5459 & T1543;
  assign T1543 = 7'h20;
  assign T5459 = T1544 ? 7'h7f : 7'h0;
  assign T1544 = T1545;
  assign T1545 = 1'h1;
  assign T5460 = T5461 ? 10'h3ff : 10'h0;
  assign T5461 = T1542[3'h6];
  assign T1546 = T1438 & T5462;
  assign T5462 = {T5463, T1547};
  assign T1547 = ~ T1543;
  assign T5463 = T5464 ? 10'h3ff : 10'h0;
  assign T5464 = T1547[3'h6];
  assign T1548 = T1458 & T1549;
  assign T1549 = 4'ha == T1457;
  assign T1550 = T1555 | T5465;
  assign T5465 = {T5467, T1551};
  assign T1551 = T5466 & T1552;
  assign T1552 = 6'h10;
  assign T5466 = T1553 ? 6'h3f : 6'h0;
  assign T1553 = T1554;
  assign T1554 = 1'h1;
  assign T5467 = T5468 ? 11'h7ff : 11'h0;
  assign T5468 = T1551[3'h5];
  assign T1555 = T1437 & T5469;
  assign T5469 = {T5470, T1556};
  assign T1556 = ~ T1552;
  assign T5470 = T5471 ? 11'h7ff : 11'h0;
  assign T5471 = T1556[3'h5];
  assign T1557 = T1458 & T1558;
  assign T1558 = 4'hb == T1457;
  assign T1559 = T1564 | T5472;
  assign T5472 = {T5474, T1560};
  assign T1560 = T5473 & T1561;
  assign T1561 = 5'h8;
  assign T5473 = T1562 ? 5'h1f : 5'h0;
  assign T1562 = T1563;
  assign T1563 = 1'h1;
  assign T5474 = T5475 ? 12'hfff : 12'h0;
  assign T5475 = T1560[3'h4];
  assign T1564 = T1436 & T5476;
  assign T5476 = {T5477, T1565};
  assign T1565 = ~ T1561;
  assign T5477 = T5478 ? 12'hfff : 12'h0;
  assign T5478 = T1565[3'h4];
  assign T1566 = T1458 & T1567;
  assign T1567 = 4'hc == T1457;
  assign T1568 = T1573 | T5479;
  assign T5479 = {T5481, T1569};
  assign T1569 = T5480 & T1570;
  assign T1570 = 4'h4;
  assign T5480 = T1571 ? 4'hf : 4'h0;
  assign T1571 = T1572;
  assign T1572 = 1'h1;
  assign T5481 = T5482 ? 13'h1fff : 13'h0;
  assign T5482 = T1569[2'h3];
  assign T1573 = T1435 & T5483;
  assign T5483 = {T5484, T1574};
  assign T1574 = ~ T1570;
  assign T5484 = T5485 ? 13'h1fff : 13'h0;
  assign T5485 = T1574[2'h3];
  assign T1575 = T1458 & T1576;
  assign T1576 = 4'hd == T1457;
  assign T1577 = T1582 | T5486;
  assign T5486 = {T5488, T1578};
  assign T1578 = T5487 & T1579;
  assign T1579 = 3'h2;
  assign T5487 = T1580 ? 3'h7 : 3'h0;
  assign T1580 = T1581;
  assign T1581 = 1'h1;
  assign T5488 = T5489 ? 14'h3fff : 14'h0;
  assign T5489 = T1578[2'h2];
  assign T1582 = T1434 & T5490;
  assign T5490 = {T5491, T1583};
  assign T1583 = ~ T1579;
  assign T5491 = T5492 ? 14'h3fff : 14'h0;
  assign T5492 = T1583[2'h2];
  assign T1584 = T1458 & T1585;
  assign T1585 = 4'he == T1457;
  assign T1586 = T1591 | T5493;
  assign T5493 = {T5495, T1587};
  assign T1587 = T5494 & T1588;
  assign T1588 = 2'h1;
  assign T5494 = T1589 ? 2'h3 : 2'h0;
  assign T1589 = T1590;
  assign T1590 = 1'h1;
  assign T5495 = T5496 ? 15'h7fff : 15'h0;
  assign T5496 = T1587[1'h1];
  assign T1591 = T1433 & T5497;
  assign T5497 = {T5498, T1592};
  assign T1592 = ~ T1588;
  assign T5498 = T5499 ? 15'h7fff : 15'h0;
  assign T5499 = T1592[1'h1];
  assign T1593 = T1458 & T1594;
  assign T1594 = 4'hf == T1457;
  assign io_V_wire_en_2 = V_wire_en_2;
  assign V_wire_en_2 = T5500;
  assign T5500 = T1595[4'hf:1'h0];
  assign T1595 = T1756 ? T1749 : T1596;
  assign T1596 = T1747 ? T1740 : T1597;
  assign T1597 = T1738 ? T1731 : T1598;
  assign T1598 = T1729 ? T1722 : T1599;
  assign T1599 = T1720 ? T1713 : T1600;
  assign T1600 = T1711 ? T1704 : T1601;
  assign T1601 = T1702 ? T1695 : T1602;
  assign T1602 = T1693 ? T1686 : T1603;
  assign T1603 = T1684 ? T1677 : T1604;
  assign T1604 = T1675 ? T1668 : T1605;
  assign T1605 = T1666 ? T1659 : T1606;
  assign T1606 = T1657 ? T1650 : T1607;
  assign T1607 = T1648 ? T1641 : T1608;
  assign T1608 = T1639 ? T1632 : T1609;
  assign T1609 = T1630 ? T1623 : T1610;
  assign T1610 = T1618 ? T1611 : 17'h0;
  assign T1611 = T1616 | T1612;
  assign T1612 = T5501 & T1613;
  assign T1613 = 17'h8000;
  assign T5501 = T1614 ? 17'h1ffff : 17'h0;
  assign T1614 = T1615;
  assign T1615 = 1'h1;
  assign T1616 = 17'h0 & T1617;
  assign T1617 = ~ T1613;
  assign T1618 = T1621 & T1619;
  assign T1619 = 4'h0 == T1620;
  assign T1620 = LogicBlockModule_2_io_config_V_out[2'h3:1'h0];
  assign T1621 = T1622;
  assign T1622 = LogicBlockModule_2_io_config_V_out[3'h4];
  assign T1623 = T1628 | T5502;
  assign T5502 = {T5504, T1624};
  assign T1624 = T5503 & T1625;
  assign T1625 = 16'h4000;
  assign T5503 = T1626 ? 16'hffff : 16'h0;
  assign T1626 = T1627;
  assign T1627 = 1'h1;
  assign T5504 = T1624[4'hf];
  assign T1628 = T1610 & T5505;
  assign T5505 = {T5506, T1629};
  assign T1629 = ~ T1625;
  assign T5506 = T1629[4'hf];
  assign T1630 = T1621 & T1631;
  assign T1631 = 4'h1 == T1620;
  assign T1632 = T1637 | T5507;
  assign T5507 = {T5509, T1633};
  assign T1633 = T5508 & T1634;
  assign T1634 = 15'h2000;
  assign T5508 = T1635 ? 15'h7fff : 15'h0;
  assign T1635 = T1636;
  assign T1636 = 1'h1;
  assign T5509 = T5510 ? 2'h3 : 2'h0;
  assign T5510 = T1633[4'he];
  assign T1637 = T1609 & T5511;
  assign T5511 = {T5512, T1638};
  assign T1638 = ~ T1634;
  assign T5512 = T5513 ? 2'h3 : 2'h0;
  assign T5513 = T1638[4'he];
  assign T1639 = T1621 & T1640;
  assign T1640 = 4'h2 == T1620;
  assign T1641 = T1646 | T5514;
  assign T5514 = {T5516, T1642};
  assign T1642 = T5515 & T1643;
  assign T1643 = 14'h1000;
  assign T5515 = T1644 ? 14'h3fff : 14'h0;
  assign T1644 = T1645;
  assign T1645 = 1'h1;
  assign T5516 = T5517 ? 3'h7 : 3'h0;
  assign T5517 = T1642[4'hd];
  assign T1646 = T1608 & T5518;
  assign T5518 = {T5519, T1647};
  assign T1647 = ~ T1643;
  assign T5519 = T5520 ? 3'h7 : 3'h0;
  assign T5520 = T1647[4'hd];
  assign T1648 = T1621 & T1649;
  assign T1649 = 4'h3 == T1620;
  assign T1650 = T1655 | T5521;
  assign T5521 = {T5523, T1651};
  assign T1651 = T5522 & T1652;
  assign T1652 = 13'h800;
  assign T5522 = T1653 ? 13'h1fff : 13'h0;
  assign T1653 = T1654;
  assign T1654 = 1'h1;
  assign T5523 = T5524 ? 4'hf : 4'h0;
  assign T5524 = T1651[4'hc];
  assign T1655 = T1607 & T5525;
  assign T5525 = {T5526, T1656};
  assign T1656 = ~ T1652;
  assign T5526 = T5527 ? 4'hf : 4'h0;
  assign T5527 = T1656[4'hc];
  assign T1657 = T1621 & T1658;
  assign T1658 = 4'h4 == T1620;
  assign T1659 = T1664 | T5528;
  assign T5528 = {T5530, T1660};
  assign T1660 = T5529 & T1661;
  assign T1661 = 12'h400;
  assign T5529 = T1662 ? 12'hfff : 12'h0;
  assign T1662 = T1663;
  assign T1663 = 1'h1;
  assign T5530 = T5531 ? 5'h1f : 5'h0;
  assign T5531 = T1660[4'hb];
  assign T1664 = T1606 & T5532;
  assign T5532 = {T5533, T1665};
  assign T1665 = ~ T1661;
  assign T5533 = T5534 ? 5'h1f : 5'h0;
  assign T5534 = T1665[4'hb];
  assign T1666 = T1621 & T1667;
  assign T1667 = 4'h5 == T1620;
  assign T1668 = T1673 | T5535;
  assign T5535 = {T5537, T1669};
  assign T1669 = T5536 & T1670;
  assign T1670 = 11'h200;
  assign T5536 = T1671 ? 11'h7ff : 11'h0;
  assign T1671 = T1672;
  assign T1672 = 1'h1;
  assign T5537 = T5538 ? 6'h3f : 6'h0;
  assign T5538 = T1669[4'ha];
  assign T1673 = T1605 & T5539;
  assign T5539 = {T5540, T1674};
  assign T1674 = ~ T1670;
  assign T5540 = T5541 ? 6'h3f : 6'h0;
  assign T5541 = T1674[4'ha];
  assign T1675 = T1621 & T1676;
  assign T1676 = 4'h6 == T1620;
  assign T1677 = T1682 | T5542;
  assign T5542 = {T5544, T1678};
  assign T1678 = T5543 & T1679;
  assign T1679 = 10'h100;
  assign T5543 = T1680 ? 10'h3ff : 10'h0;
  assign T1680 = T1681;
  assign T1681 = 1'h1;
  assign T5544 = T5545 ? 7'h7f : 7'h0;
  assign T5545 = T1678[4'h9];
  assign T1682 = T1604 & T5546;
  assign T5546 = {T5547, T1683};
  assign T1683 = ~ T1679;
  assign T5547 = T5548 ? 7'h7f : 7'h0;
  assign T5548 = T1683[4'h9];
  assign T1684 = T1621 & T1685;
  assign T1685 = 4'h7 == T1620;
  assign T1686 = T1691 | T5549;
  assign T5549 = {T5551, T1687};
  assign T1687 = T5550 & T1688;
  assign T1688 = 9'h80;
  assign T5550 = T1689 ? 9'h1ff : 9'h0;
  assign T1689 = T1690;
  assign T1690 = 1'h1;
  assign T5551 = T5552 ? 8'hff : 8'h0;
  assign T5552 = T1687[4'h8];
  assign T1691 = T1603 & T5553;
  assign T5553 = {T5554, T1692};
  assign T1692 = ~ T1688;
  assign T5554 = T5555 ? 8'hff : 8'h0;
  assign T5555 = T1692[4'h8];
  assign T1693 = T1621 & T1694;
  assign T1694 = 4'h8 == T1620;
  assign T1695 = T1700 | T5556;
  assign T5556 = {T5558, T1696};
  assign T1696 = T5557 & T1697;
  assign T1697 = 8'h40;
  assign T5557 = T1698 ? 8'hff : 8'h0;
  assign T1698 = T1699;
  assign T1699 = 1'h1;
  assign T5558 = T5559 ? 9'h1ff : 9'h0;
  assign T5559 = T1696[3'h7];
  assign T1700 = T1602 & T5560;
  assign T5560 = {T5561, T1701};
  assign T1701 = ~ T1697;
  assign T5561 = T5562 ? 9'h1ff : 9'h0;
  assign T5562 = T1701[3'h7];
  assign T1702 = T1621 & T1703;
  assign T1703 = 4'h9 == T1620;
  assign T1704 = T1709 | T5563;
  assign T5563 = {T5565, T1705};
  assign T1705 = T5564 & T1706;
  assign T1706 = 7'h20;
  assign T5564 = T1707 ? 7'h7f : 7'h0;
  assign T1707 = T1708;
  assign T1708 = 1'h1;
  assign T5565 = T5566 ? 10'h3ff : 10'h0;
  assign T5566 = T1705[3'h6];
  assign T1709 = T1601 & T5567;
  assign T5567 = {T5568, T1710};
  assign T1710 = ~ T1706;
  assign T5568 = T5569 ? 10'h3ff : 10'h0;
  assign T5569 = T1710[3'h6];
  assign T1711 = T1621 & T1712;
  assign T1712 = 4'ha == T1620;
  assign T1713 = T1718 | T5570;
  assign T5570 = {T5572, T1714};
  assign T1714 = T5571 & T1715;
  assign T1715 = 6'h10;
  assign T5571 = T1716 ? 6'h3f : 6'h0;
  assign T1716 = T1717;
  assign T1717 = 1'h1;
  assign T5572 = T5573 ? 11'h7ff : 11'h0;
  assign T5573 = T1714[3'h5];
  assign T1718 = T1600 & T5574;
  assign T5574 = {T5575, T1719};
  assign T1719 = ~ T1715;
  assign T5575 = T5576 ? 11'h7ff : 11'h0;
  assign T5576 = T1719[3'h5];
  assign T1720 = T1621 & T1721;
  assign T1721 = 4'hb == T1620;
  assign T1722 = T1727 | T5577;
  assign T5577 = {T5579, T1723};
  assign T1723 = T5578 & T1724;
  assign T1724 = 5'h8;
  assign T5578 = T1725 ? 5'h1f : 5'h0;
  assign T1725 = T1726;
  assign T1726 = 1'h1;
  assign T5579 = T5580 ? 12'hfff : 12'h0;
  assign T5580 = T1723[3'h4];
  assign T1727 = T1599 & T5581;
  assign T5581 = {T5582, T1728};
  assign T1728 = ~ T1724;
  assign T5582 = T5583 ? 12'hfff : 12'h0;
  assign T5583 = T1728[3'h4];
  assign T1729 = T1621 & T1730;
  assign T1730 = 4'hc == T1620;
  assign T1731 = T1736 | T5584;
  assign T5584 = {T5586, T1732};
  assign T1732 = T5585 & T1733;
  assign T1733 = 4'h4;
  assign T5585 = T1734 ? 4'hf : 4'h0;
  assign T1734 = T1735;
  assign T1735 = 1'h1;
  assign T5586 = T5587 ? 13'h1fff : 13'h0;
  assign T5587 = T1732[2'h3];
  assign T1736 = T1598 & T5588;
  assign T5588 = {T5589, T1737};
  assign T1737 = ~ T1733;
  assign T5589 = T5590 ? 13'h1fff : 13'h0;
  assign T5590 = T1737[2'h3];
  assign T1738 = T1621 & T1739;
  assign T1739 = 4'hd == T1620;
  assign T1740 = T1745 | T5591;
  assign T5591 = {T5593, T1741};
  assign T1741 = T5592 & T1742;
  assign T1742 = 3'h2;
  assign T5592 = T1743 ? 3'h7 : 3'h0;
  assign T1743 = T1744;
  assign T1744 = 1'h1;
  assign T5593 = T5594 ? 14'h3fff : 14'h0;
  assign T5594 = T1741[2'h2];
  assign T1745 = T1597 & T5595;
  assign T5595 = {T5596, T1746};
  assign T1746 = ~ T1742;
  assign T5596 = T5597 ? 14'h3fff : 14'h0;
  assign T5597 = T1746[2'h2];
  assign T1747 = T1621 & T1748;
  assign T1748 = 4'he == T1620;
  assign T1749 = T1754 | T5598;
  assign T5598 = {T5600, T1750};
  assign T1750 = T5599 & T1751;
  assign T1751 = 2'h1;
  assign T5599 = T1752 ? 2'h3 : 2'h0;
  assign T1752 = T1753;
  assign T1753 = 1'h1;
  assign T5600 = T5601 ? 15'h7fff : 15'h0;
  assign T5601 = T1750[1'h1];
  assign T1754 = T1596 & T5602;
  assign T5602 = {T5603, T1755};
  assign T1755 = ~ T1751;
  assign T5603 = T5604 ? 15'h7fff : 15'h0;
  assign T5604 = T1755[1'h1];
  assign T1756 = T1621 & T1757;
  assign T1757 = 4'hf == T1620;
  assign io_V_wire_en_3 = V_wire_en_3;
  assign V_wire_en_3 = T5605;
  assign T5605 = T1758[4'hf:1'h0];
  assign T1758 = T1919 ? T1912 : T1759;
  assign T1759 = T1910 ? T1903 : T1760;
  assign T1760 = T1901 ? T1894 : T1761;
  assign T1761 = T1892 ? T1885 : T1762;
  assign T1762 = T1883 ? T1876 : T1763;
  assign T1763 = T1874 ? T1867 : T1764;
  assign T1764 = T1865 ? T1858 : T1765;
  assign T1765 = T1856 ? T1849 : T1766;
  assign T1766 = T1847 ? T1840 : T1767;
  assign T1767 = T1838 ? T1831 : T1768;
  assign T1768 = T1829 ? T1822 : T1769;
  assign T1769 = T1820 ? T1813 : T1770;
  assign T1770 = T1811 ? T1804 : T1771;
  assign T1771 = T1802 ? T1795 : T1772;
  assign T1772 = T1793 ? T1786 : T1773;
  assign T1773 = T1781 ? T1774 : 17'h0;
  assign T1774 = T1779 | T1775;
  assign T1775 = T5606 & T1776;
  assign T1776 = 17'h8000;
  assign T5606 = T1777 ? 17'h1ffff : 17'h0;
  assign T1777 = T1778;
  assign T1778 = 1'h1;
  assign T1779 = 17'h0 & T1780;
  assign T1780 = ~ T1776;
  assign T1781 = T1784 & T1782;
  assign T1782 = 4'h0 == T1783;
  assign T1783 = LogicBlockModule_3_io_config_V_out[2'h3:1'h0];
  assign T1784 = T1785;
  assign T1785 = LogicBlockModule_3_io_config_V_out[3'h4];
  assign T1786 = T1791 | T5607;
  assign T5607 = {T5609, T1787};
  assign T1787 = T5608 & T1788;
  assign T1788 = 16'h4000;
  assign T5608 = T1789 ? 16'hffff : 16'h0;
  assign T1789 = T1790;
  assign T1790 = 1'h1;
  assign T5609 = T1787[4'hf];
  assign T1791 = T1773 & T5610;
  assign T5610 = {T5611, T1792};
  assign T1792 = ~ T1788;
  assign T5611 = T1792[4'hf];
  assign T1793 = T1784 & T1794;
  assign T1794 = 4'h1 == T1783;
  assign T1795 = T1800 | T5612;
  assign T5612 = {T5614, T1796};
  assign T1796 = T5613 & T1797;
  assign T1797 = 15'h2000;
  assign T5613 = T1798 ? 15'h7fff : 15'h0;
  assign T1798 = T1799;
  assign T1799 = 1'h1;
  assign T5614 = T5615 ? 2'h3 : 2'h0;
  assign T5615 = T1796[4'he];
  assign T1800 = T1772 & T5616;
  assign T5616 = {T5617, T1801};
  assign T1801 = ~ T1797;
  assign T5617 = T5618 ? 2'h3 : 2'h0;
  assign T5618 = T1801[4'he];
  assign T1802 = T1784 & T1803;
  assign T1803 = 4'h2 == T1783;
  assign T1804 = T1809 | T5619;
  assign T5619 = {T5621, T1805};
  assign T1805 = T5620 & T1806;
  assign T1806 = 14'h1000;
  assign T5620 = T1807 ? 14'h3fff : 14'h0;
  assign T1807 = T1808;
  assign T1808 = 1'h1;
  assign T5621 = T5622 ? 3'h7 : 3'h0;
  assign T5622 = T1805[4'hd];
  assign T1809 = T1771 & T5623;
  assign T5623 = {T5624, T1810};
  assign T1810 = ~ T1806;
  assign T5624 = T5625 ? 3'h7 : 3'h0;
  assign T5625 = T1810[4'hd];
  assign T1811 = T1784 & T1812;
  assign T1812 = 4'h3 == T1783;
  assign T1813 = T1818 | T5626;
  assign T5626 = {T5628, T1814};
  assign T1814 = T5627 & T1815;
  assign T1815 = 13'h800;
  assign T5627 = T1816 ? 13'h1fff : 13'h0;
  assign T1816 = T1817;
  assign T1817 = 1'h1;
  assign T5628 = T5629 ? 4'hf : 4'h0;
  assign T5629 = T1814[4'hc];
  assign T1818 = T1770 & T5630;
  assign T5630 = {T5631, T1819};
  assign T1819 = ~ T1815;
  assign T5631 = T5632 ? 4'hf : 4'h0;
  assign T5632 = T1819[4'hc];
  assign T1820 = T1784 & T1821;
  assign T1821 = 4'h4 == T1783;
  assign T1822 = T1827 | T5633;
  assign T5633 = {T5635, T1823};
  assign T1823 = T5634 & T1824;
  assign T1824 = 12'h400;
  assign T5634 = T1825 ? 12'hfff : 12'h0;
  assign T1825 = T1826;
  assign T1826 = 1'h1;
  assign T5635 = T5636 ? 5'h1f : 5'h0;
  assign T5636 = T1823[4'hb];
  assign T1827 = T1769 & T5637;
  assign T5637 = {T5638, T1828};
  assign T1828 = ~ T1824;
  assign T5638 = T5639 ? 5'h1f : 5'h0;
  assign T5639 = T1828[4'hb];
  assign T1829 = T1784 & T1830;
  assign T1830 = 4'h5 == T1783;
  assign T1831 = T1836 | T5640;
  assign T5640 = {T5642, T1832};
  assign T1832 = T5641 & T1833;
  assign T1833 = 11'h200;
  assign T5641 = T1834 ? 11'h7ff : 11'h0;
  assign T1834 = T1835;
  assign T1835 = 1'h1;
  assign T5642 = T5643 ? 6'h3f : 6'h0;
  assign T5643 = T1832[4'ha];
  assign T1836 = T1768 & T5644;
  assign T5644 = {T5645, T1837};
  assign T1837 = ~ T1833;
  assign T5645 = T5646 ? 6'h3f : 6'h0;
  assign T5646 = T1837[4'ha];
  assign T1838 = T1784 & T1839;
  assign T1839 = 4'h6 == T1783;
  assign T1840 = T1845 | T5647;
  assign T5647 = {T5649, T1841};
  assign T1841 = T5648 & T1842;
  assign T1842 = 10'h100;
  assign T5648 = T1843 ? 10'h3ff : 10'h0;
  assign T1843 = T1844;
  assign T1844 = 1'h1;
  assign T5649 = T5650 ? 7'h7f : 7'h0;
  assign T5650 = T1841[4'h9];
  assign T1845 = T1767 & T5651;
  assign T5651 = {T5652, T1846};
  assign T1846 = ~ T1842;
  assign T5652 = T5653 ? 7'h7f : 7'h0;
  assign T5653 = T1846[4'h9];
  assign T1847 = T1784 & T1848;
  assign T1848 = 4'h7 == T1783;
  assign T1849 = T1854 | T5654;
  assign T5654 = {T5656, T1850};
  assign T1850 = T5655 & T1851;
  assign T1851 = 9'h80;
  assign T5655 = T1852 ? 9'h1ff : 9'h0;
  assign T1852 = T1853;
  assign T1853 = 1'h1;
  assign T5656 = T5657 ? 8'hff : 8'h0;
  assign T5657 = T1850[4'h8];
  assign T1854 = T1766 & T5658;
  assign T5658 = {T5659, T1855};
  assign T1855 = ~ T1851;
  assign T5659 = T5660 ? 8'hff : 8'h0;
  assign T5660 = T1855[4'h8];
  assign T1856 = T1784 & T1857;
  assign T1857 = 4'h8 == T1783;
  assign T1858 = T1863 | T5661;
  assign T5661 = {T5663, T1859};
  assign T1859 = T5662 & T1860;
  assign T1860 = 8'h40;
  assign T5662 = T1861 ? 8'hff : 8'h0;
  assign T1861 = T1862;
  assign T1862 = 1'h1;
  assign T5663 = T5664 ? 9'h1ff : 9'h0;
  assign T5664 = T1859[3'h7];
  assign T1863 = T1765 & T5665;
  assign T5665 = {T5666, T1864};
  assign T1864 = ~ T1860;
  assign T5666 = T5667 ? 9'h1ff : 9'h0;
  assign T5667 = T1864[3'h7];
  assign T1865 = T1784 & T1866;
  assign T1866 = 4'h9 == T1783;
  assign T1867 = T1872 | T5668;
  assign T5668 = {T5670, T1868};
  assign T1868 = T5669 & T1869;
  assign T1869 = 7'h20;
  assign T5669 = T1870 ? 7'h7f : 7'h0;
  assign T1870 = T1871;
  assign T1871 = 1'h1;
  assign T5670 = T5671 ? 10'h3ff : 10'h0;
  assign T5671 = T1868[3'h6];
  assign T1872 = T1764 & T5672;
  assign T5672 = {T5673, T1873};
  assign T1873 = ~ T1869;
  assign T5673 = T5674 ? 10'h3ff : 10'h0;
  assign T5674 = T1873[3'h6];
  assign T1874 = T1784 & T1875;
  assign T1875 = 4'ha == T1783;
  assign T1876 = T1881 | T5675;
  assign T5675 = {T5677, T1877};
  assign T1877 = T5676 & T1878;
  assign T1878 = 6'h10;
  assign T5676 = T1879 ? 6'h3f : 6'h0;
  assign T1879 = T1880;
  assign T1880 = 1'h1;
  assign T5677 = T5678 ? 11'h7ff : 11'h0;
  assign T5678 = T1877[3'h5];
  assign T1881 = T1763 & T5679;
  assign T5679 = {T5680, T1882};
  assign T1882 = ~ T1878;
  assign T5680 = T5681 ? 11'h7ff : 11'h0;
  assign T5681 = T1882[3'h5];
  assign T1883 = T1784 & T1884;
  assign T1884 = 4'hb == T1783;
  assign T1885 = T1890 | T5682;
  assign T5682 = {T5684, T1886};
  assign T1886 = T5683 & T1887;
  assign T1887 = 5'h8;
  assign T5683 = T1888 ? 5'h1f : 5'h0;
  assign T1888 = T1889;
  assign T1889 = 1'h1;
  assign T5684 = T5685 ? 12'hfff : 12'h0;
  assign T5685 = T1886[3'h4];
  assign T1890 = T1762 & T5686;
  assign T5686 = {T5687, T1891};
  assign T1891 = ~ T1887;
  assign T5687 = T5688 ? 12'hfff : 12'h0;
  assign T5688 = T1891[3'h4];
  assign T1892 = T1784 & T1893;
  assign T1893 = 4'hc == T1783;
  assign T1894 = T1899 | T5689;
  assign T5689 = {T5691, T1895};
  assign T1895 = T5690 & T1896;
  assign T1896 = 4'h4;
  assign T5690 = T1897 ? 4'hf : 4'h0;
  assign T1897 = T1898;
  assign T1898 = 1'h1;
  assign T5691 = T5692 ? 13'h1fff : 13'h0;
  assign T5692 = T1895[2'h3];
  assign T1899 = T1761 & T5693;
  assign T5693 = {T5694, T1900};
  assign T1900 = ~ T1896;
  assign T5694 = T5695 ? 13'h1fff : 13'h0;
  assign T5695 = T1900[2'h3];
  assign T1901 = T1784 & T1902;
  assign T1902 = 4'hd == T1783;
  assign T1903 = T1908 | T5696;
  assign T5696 = {T5698, T1904};
  assign T1904 = T5697 & T1905;
  assign T1905 = 3'h2;
  assign T5697 = T1906 ? 3'h7 : 3'h0;
  assign T1906 = T1907;
  assign T1907 = 1'h1;
  assign T5698 = T5699 ? 14'h3fff : 14'h0;
  assign T5699 = T1904[2'h2];
  assign T1908 = T1760 & T5700;
  assign T5700 = {T5701, T1909};
  assign T1909 = ~ T1905;
  assign T5701 = T5702 ? 14'h3fff : 14'h0;
  assign T5702 = T1909[2'h2];
  assign T1910 = T1784 & T1911;
  assign T1911 = 4'he == T1783;
  assign T1912 = T1917 | T5703;
  assign T5703 = {T5705, T1913};
  assign T1913 = T5704 & T1914;
  assign T1914 = 2'h1;
  assign T5704 = T1915 ? 2'h3 : 2'h0;
  assign T1915 = T1916;
  assign T1916 = 1'h1;
  assign T5705 = T5706 ? 15'h7fff : 15'h0;
  assign T5706 = T1913[1'h1];
  assign T1917 = T1759 & T5707;
  assign T5707 = {T5708, T1918};
  assign T1918 = ~ T1914;
  assign T5708 = T5709 ? 15'h7fff : 15'h0;
  assign T5709 = T1918[1'h1];
  assign T1919 = T1784 & T1920;
  assign T1920 = 4'hf == T1783;
  assign io_V_wire_en_4 = V_wire_en_4;
  assign V_wire_en_4 = T5710;
  assign T5710 = T1921[4'hf:1'h0];
  assign T1921 = T2082 ? T2075 : T1922;
  assign T1922 = T2073 ? T2066 : T1923;
  assign T1923 = T2064 ? T2057 : T1924;
  assign T1924 = T2055 ? T2048 : T1925;
  assign T1925 = T2046 ? T2039 : T1926;
  assign T1926 = T2037 ? T2030 : T1927;
  assign T1927 = T2028 ? T2021 : T1928;
  assign T1928 = T2019 ? T2012 : T1929;
  assign T1929 = T2010 ? T2003 : T1930;
  assign T1930 = T2001 ? T1994 : T1931;
  assign T1931 = T1992 ? T1985 : T1932;
  assign T1932 = T1983 ? T1976 : T1933;
  assign T1933 = T1974 ? T1967 : T1934;
  assign T1934 = T1965 ? T1958 : T1935;
  assign T1935 = T1956 ? T1949 : T1936;
  assign T1936 = T1944 ? T1937 : 17'h0;
  assign T1937 = T1942 | T1938;
  assign T1938 = T5711 & T1939;
  assign T1939 = 17'h8000;
  assign T5711 = T1940 ? 17'h1ffff : 17'h0;
  assign T1940 = T1941;
  assign T1941 = 1'h1;
  assign T1942 = 17'h0 & T1943;
  assign T1943 = ~ T1939;
  assign T1944 = T1947 & T1945;
  assign T1945 = 4'h0 == T1946;
  assign T1946 = LogicBlockModule_4_io_config_V_out[2'h3:1'h0];
  assign T1947 = T1948;
  assign T1948 = LogicBlockModule_4_io_config_V_out[3'h4];
  assign T1949 = T1954 | T5712;
  assign T5712 = {T5714, T1950};
  assign T1950 = T5713 & T1951;
  assign T1951 = 16'h4000;
  assign T5713 = T1952 ? 16'hffff : 16'h0;
  assign T1952 = T1953;
  assign T1953 = 1'h1;
  assign T5714 = T1950[4'hf];
  assign T1954 = T1936 & T5715;
  assign T5715 = {T5716, T1955};
  assign T1955 = ~ T1951;
  assign T5716 = T1955[4'hf];
  assign T1956 = T1947 & T1957;
  assign T1957 = 4'h1 == T1946;
  assign T1958 = T1963 | T5717;
  assign T5717 = {T5719, T1959};
  assign T1959 = T5718 & T1960;
  assign T1960 = 15'h2000;
  assign T5718 = T1961 ? 15'h7fff : 15'h0;
  assign T1961 = T1962;
  assign T1962 = 1'h1;
  assign T5719 = T5720 ? 2'h3 : 2'h0;
  assign T5720 = T1959[4'he];
  assign T1963 = T1935 & T5721;
  assign T5721 = {T5722, T1964};
  assign T1964 = ~ T1960;
  assign T5722 = T5723 ? 2'h3 : 2'h0;
  assign T5723 = T1964[4'he];
  assign T1965 = T1947 & T1966;
  assign T1966 = 4'h2 == T1946;
  assign T1967 = T1972 | T5724;
  assign T5724 = {T5726, T1968};
  assign T1968 = T5725 & T1969;
  assign T1969 = 14'h1000;
  assign T5725 = T1970 ? 14'h3fff : 14'h0;
  assign T1970 = T1971;
  assign T1971 = 1'h1;
  assign T5726 = T5727 ? 3'h7 : 3'h0;
  assign T5727 = T1968[4'hd];
  assign T1972 = T1934 & T5728;
  assign T5728 = {T5729, T1973};
  assign T1973 = ~ T1969;
  assign T5729 = T5730 ? 3'h7 : 3'h0;
  assign T5730 = T1973[4'hd];
  assign T1974 = T1947 & T1975;
  assign T1975 = 4'h3 == T1946;
  assign T1976 = T1981 | T5731;
  assign T5731 = {T5733, T1977};
  assign T1977 = T5732 & T1978;
  assign T1978 = 13'h800;
  assign T5732 = T1979 ? 13'h1fff : 13'h0;
  assign T1979 = T1980;
  assign T1980 = 1'h1;
  assign T5733 = T5734 ? 4'hf : 4'h0;
  assign T5734 = T1977[4'hc];
  assign T1981 = T1933 & T5735;
  assign T5735 = {T5736, T1982};
  assign T1982 = ~ T1978;
  assign T5736 = T5737 ? 4'hf : 4'h0;
  assign T5737 = T1982[4'hc];
  assign T1983 = T1947 & T1984;
  assign T1984 = 4'h4 == T1946;
  assign T1985 = T1990 | T5738;
  assign T5738 = {T5740, T1986};
  assign T1986 = T5739 & T1987;
  assign T1987 = 12'h400;
  assign T5739 = T1988 ? 12'hfff : 12'h0;
  assign T1988 = T1989;
  assign T1989 = 1'h1;
  assign T5740 = T5741 ? 5'h1f : 5'h0;
  assign T5741 = T1986[4'hb];
  assign T1990 = T1932 & T5742;
  assign T5742 = {T5743, T1991};
  assign T1991 = ~ T1987;
  assign T5743 = T5744 ? 5'h1f : 5'h0;
  assign T5744 = T1991[4'hb];
  assign T1992 = T1947 & T1993;
  assign T1993 = 4'h5 == T1946;
  assign T1994 = T1999 | T5745;
  assign T5745 = {T5747, T1995};
  assign T1995 = T5746 & T1996;
  assign T1996 = 11'h200;
  assign T5746 = T1997 ? 11'h7ff : 11'h0;
  assign T1997 = T1998;
  assign T1998 = 1'h1;
  assign T5747 = T5748 ? 6'h3f : 6'h0;
  assign T5748 = T1995[4'ha];
  assign T1999 = T1931 & T5749;
  assign T5749 = {T5750, T2000};
  assign T2000 = ~ T1996;
  assign T5750 = T5751 ? 6'h3f : 6'h0;
  assign T5751 = T2000[4'ha];
  assign T2001 = T1947 & T2002;
  assign T2002 = 4'h6 == T1946;
  assign T2003 = T2008 | T5752;
  assign T5752 = {T5754, T2004};
  assign T2004 = T5753 & T2005;
  assign T2005 = 10'h100;
  assign T5753 = T2006 ? 10'h3ff : 10'h0;
  assign T2006 = T2007;
  assign T2007 = 1'h1;
  assign T5754 = T5755 ? 7'h7f : 7'h0;
  assign T5755 = T2004[4'h9];
  assign T2008 = T1930 & T5756;
  assign T5756 = {T5757, T2009};
  assign T2009 = ~ T2005;
  assign T5757 = T5758 ? 7'h7f : 7'h0;
  assign T5758 = T2009[4'h9];
  assign T2010 = T1947 & T2011;
  assign T2011 = 4'h7 == T1946;
  assign T2012 = T2017 | T5759;
  assign T5759 = {T5761, T2013};
  assign T2013 = T5760 & T2014;
  assign T2014 = 9'h80;
  assign T5760 = T2015 ? 9'h1ff : 9'h0;
  assign T2015 = T2016;
  assign T2016 = 1'h1;
  assign T5761 = T5762 ? 8'hff : 8'h0;
  assign T5762 = T2013[4'h8];
  assign T2017 = T1929 & T5763;
  assign T5763 = {T5764, T2018};
  assign T2018 = ~ T2014;
  assign T5764 = T5765 ? 8'hff : 8'h0;
  assign T5765 = T2018[4'h8];
  assign T2019 = T1947 & T2020;
  assign T2020 = 4'h8 == T1946;
  assign T2021 = T2026 | T5766;
  assign T5766 = {T5768, T2022};
  assign T2022 = T5767 & T2023;
  assign T2023 = 8'h40;
  assign T5767 = T2024 ? 8'hff : 8'h0;
  assign T2024 = T2025;
  assign T2025 = 1'h1;
  assign T5768 = T5769 ? 9'h1ff : 9'h0;
  assign T5769 = T2022[3'h7];
  assign T2026 = T1928 & T5770;
  assign T5770 = {T5771, T2027};
  assign T2027 = ~ T2023;
  assign T5771 = T5772 ? 9'h1ff : 9'h0;
  assign T5772 = T2027[3'h7];
  assign T2028 = T1947 & T2029;
  assign T2029 = 4'h9 == T1946;
  assign T2030 = T2035 | T5773;
  assign T5773 = {T5775, T2031};
  assign T2031 = T5774 & T2032;
  assign T2032 = 7'h20;
  assign T5774 = T2033 ? 7'h7f : 7'h0;
  assign T2033 = T2034;
  assign T2034 = 1'h1;
  assign T5775 = T5776 ? 10'h3ff : 10'h0;
  assign T5776 = T2031[3'h6];
  assign T2035 = T1927 & T5777;
  assign T5777 = {T5778, T2036};
  assign T2036 = ~ T2032;
  assign T5778 = T5779 ? 10'h3ff : 10'h0;
  assign T5779 = T2036[3'h6];
  assign T2037 = T1947 & T2038;
  assign T2038 = 4'ha == T1946;
  assign T2039 = T2044 | T5780;
  assign T5780 = {T5782, T2040};
  assign T2040 = T5781 & T2041;
  assign T2041 = 6'h10;
  assign T5781 = T2042 ? 6'h3f : 6'h0;
  assign T2042 = T2043;
  assign T2043 = 1'h1;
  assign T5782 = T5783 ? 11'h7ff : 11'h0;
  assign T5783 = T2040[3'h5];
  assign T2044 = T1926 & T5784;
  assign T5784 = {T5785, T2045};
  assign T2045 = ~ T2041;
  assign T5785 = T5786 ? 11'h7ff : 11'h0;
  assign T5786 = T2045[3'h5];
  assign T2046 = T1947 & T2047;
  assign T2047 = 4'hb == T1946;
  assign T2048 = T2053 | T5787;
  assign T5787 = {T5789, T2049};
  assign T2049 = T5788 & T2050;
  assign T2050 = 5'h8;
  assign T5788 = T2051 ? 5'h1f : 5'h0;
  assign T2051 = T2052;
  assign T2052 = 1'h1;
  assign T5789 = T5790 ? 12'hfff : 12'h0;
  assign T5790 = T2049[3'h4];
  assign T2053 = T1925 & T5791;
  assign T5791 = {T5792, T2054};
  assign T2054 = ~ T2050;
  assign T5792 = T5793 ? 12'hfff : 12'h0;
  assign T5793 = T2054[3'h4];
  assign T2055 = T1947 & T2056;
  assign T2056 = 4'hc == T1946;
  assign T2057 = T2062 | T5794;
  assign T5794 = {T5796, T2058};
  assign T2058 = T5795 & T2059;
  assign T2059 = 4'h4;
  assign T5795 = T2060 ? 4'hf : 4'h0;
  assign T2060 = T2061;
  assign T2061 = 1'h1;
  assign T5796 = T5797 ? 13'h1fff : 13'h0;
  assign T5797 = T2058[2'h3];
  assign T2062 = T1924 & T5798;
  assign T5798 = {T5799, T2063};
  assign T2063 = ~ T2059;
  assign T5799 = T5800 ? 13'h1fff : 13'h0;
  assign T5800 = T2063[2'h3];
  assign T2064 = T1947 & T2065;
  assign T2065 = 4'hd == T1946;
  assign T2066 = T2071 | T5801;
  assign T5801 = {T5803, T2067};
  assign T2067 = T5802 & T2068;
  assign T2068 = 3'h2;
  assign T5802 = T2069 ? 3'h7 : 3'h0;
  assign T2069 = T2070;
  assign T2070 = 1'h1;
  assign T5803 = T5804 ? 14'h3fff : 14'h0;
  assign T5804 = T2067[2'h2];
  assign T2071 = T1923 & T5805;
  assign T5805 = {T5806, T2072};
  assign T2072 = ~ T2068;
  assign T5806 = T5807 ? 14'h3fff : 14'h0;
  assign T5807 = T2072[2'h2];
  assign T2073 = T1947 & T2074;
  assign T2074 = 4'he == T1946;
  assign T2075 = T2080 | T5808;
  assign T5808 = {T5810, T2076};
  assign T2076 = T5809 & T2077;
  assign T2077 = 2'h1;
  assign T5809 = T2078 ? 2'h3 : 2'h0;
  assign T2078 = T2079;
  assign T2079 = 1'h1;
  assign T5810 = T5811 ? 15'h7fff : 15'h0;
  assign T5811 = T2076[1'h1];
  assign T2080 = T1922 & T5812;
  assign T5812 = {T5813, T2081};
  assign T2081 = ~ T2077;
  assign T5813 = T5814 ? 15'h7fff : 15'h0;
  assign T5814 = T2081[1'h1];
  assign T2082 = T1947 & T2083;
  assign T2083 = 4'hf == T1946;
  assign io_V_wire_en_5 = V_wire_en_5;
  assign V_wire_en_5 = T5815;
  assign T5815 = T2084[4'hf:1'h0];
  assign T2084 = T2245 ? T2238 : T2085;
  assign T2085 = T2236 ? T2229 : T2086;
  assign T2086 = T2227 ? T2220 : T2087;
  assign T2087 = T2218 ? T2211 : T2088;
  assign T2088 = T2209 ? T2202 : T2089;
  assign T2089 = T2200 ? T2193 : T2090;
  assign T2090 = T2191 ? T2184 : T2091;
  assign T2091 = T2182 ? T2175 : T2092;
  assign T2092 = T2173 ? T2166 : T2093;
  assign T2093 = T2164 ? T2157 : T2094;
  assign T2094 = T2155 ? T2148 : T2095;
  assign T2095 = T2146 ? T2139 : T2096;
  assign T2096 = T2137 ? T2130 : T2097;
  assign T2097 = T2128 ? T2121 : T2098;
  assign T2098 = T2119 ? T2112 : T2099;
  assign T2099 = T2107 ? T2100 : 17'h0;
  assign T2100 = T2105 | T2101;
  assign T2101 = T5816 & T2102;
  assign T2102 = 17'h8000;
  assign T5816 = T2103 ? 17'h1ffff : 17'h0;
  assign T2103 = T2104;
  assign T2104 = 1'h1;
  assign T2105 = 17'h0 & T2106;
  assign T2106 = ~ T2102;
  assign T2107 = T2110 & T2108;
  assign T2108 = 4'h0 == T2109;
  assign T2109 = LogicBlockModule_5_io_config_V_out[2'h3:1'h0];
  assign T2110 = T2111;
  assign T2111 = LogicBlockModule_5_io_config_V_out[3'h4];
  assign T2112 = T2117 | T5817;
  assign T5817 = {T5819, T2113};
  assign T2113 = T5818 & T2114;
  assign T2114 = 16'h4000;
  assign T5818 = T2115 ? 16'hffff : 16'h0;
  assign T2115 = T2116;
  assign T2116 = 1'h1;
  assign T5819 = T2113[4'hf];
  assign T2117 = T2099 & T5820;
  assign T5820 = {T5821, T2118};
  assign T2118 = ~ T2114;
  assign T5821 = T2118[4'hf];
  assign T2119 = T2110 & T2120;
  assign T2120 = 4'h1 == T2109;
  assign T2121 = T2126 | T5822;
  assign T5822 = {T5824, T2122};
  assign T2122 = T5823 & T2123;
  assign T2123 = 15'h2000;
  assign T5823 = T2124 ? 15'h7fff : 15'h0;
  assign T2124 = T2125;
  assign T2125 = 1'h1;
  assign T5824 = T5825 ? 2'h3 : 2'h0;
  assign T5825 = T2122[4'he];
  assign T2126 = T2098 & T5826;
  assign T5826 = {T5827, T2127};
  assign T2127 = ~ T2123;
  assign T5827 = T5828 ? 2'h3 : 2'h0;
  assign T5828 = T2127[4'he];
  assign T2128 = T2110 & T2129;
  assign T2129 = 4'h2 == T2109;
  assign T2130 = T2135 | T5829;
  assign T5829 = {T5831, T2131};
  assign T2131 = T5830 & T2132;
  assign T2132 = 14'h1000;
  assign T5830 = T2133 ? 14'h3fff : 14'h0;
  assign T2133 = T2134;
  assign T2134 = 1'h1;
  assign T5831 = T5832 ? 3'h7 : 3'h0;
  assign T5832 = T2131[4'hd];
  assign T2135 = T2097 & T5833;
  assign T5833 = {T5834, T2136};
  assign T2136 = ~ T2132;
  assign T5834 = T5835 ? 3'h7 : 3'h0;
  assign T5835 = T2136[4'hd];
  assign T2137 = T2110 & T2138;
  assign T2138 = 4'h3 == T2109;
  assign T2139 = T2144 | T5836;
  assign T5836 = {T5838, T2140};
  assign T2140 = T5837 & T2141;
  assign T2141 = 13'h800;
  assign T5837 = T2142 ? 13'h1fff : 13'h0;
  assign T2142 = T2143;
  assign T2143 = 1'h1;
  assign T5838 = T5839 ? 4'hf : 4'h0;
  assign T5839 = T2140[4'hc];
  assign T2144 = T2096 & T5840;
  assign T5840 = {T5841, T2145};
  assign T2145 = ~ T2141;
  assign T5841 = T5842 ? 4'hf : 4'h0;
  assign T5842 = T2145[4'hc];
  assign T2146 = T2110 & T2147;
  assign T2147 = 4'h4 == T2109;
  assign T2148 = T2153 | T5843;
  assign T5843 = {T5845, T2149};
  assign T2149 = T5844 & T2150;
  assign T2150 = 12'h400;
  assign T5844 = T2151 ? 12'hfff : 12'h0;
  assign T2151 = T2152;
  assign T2152 = 1'h1;
  assign T5845 = T5846 ? 5'h1f : 5'h0;
  assign T5846 = T2149[4'hb];
  assign T2153 = T2095 & T5847;
  assign T5847 = {T5848, T2154};
  assign T2154 = ~ T2150;
  assign T5848 = T5849 ? 5'h1f : 5'h0;
  assign T5849 = T2154[4'hb];
  assign T2155 = T2110 & T2156;
  assign T2156 = 4'h5 == T2109;
  assign T2157 = T2162 | T5850;
  assign T5850 = {T5852, T2158};
  assign T2158 = T5851 & T2159;
  assign T2159 = 11'h200;
  assign T5851 = T2160 ? 11'h7ff : 11'h0;
  assign T2160 = T2161;
  assign T2161 = 1'h1;
  assign T5852 = T5853 ? 6'h3f : 6'h0;
  assign T5853 = T2158[4'ha];
  assign T2162 = T2094 & T5854;
  assign T5854 = {T5855, T2163};
  assign T2163 = ~ T2159;
  assign T5855 = T5856 ? 6'h3f : 6'h0;
  assign T5856 = T2163[4'ha];
  assign T2164 = T2110 & T2165;
  assign T2165 = 4'h6 == T2109;
  assign T2166 = T2171 | T5857;
  assign T5857 = {T5859, T2167};
  assign T2167 = T5858 & T2168;
  assign T2168 = 10'h100;
  assign T5858 = T2169 ? 10'h3ff : 10'h0;
  assign T2169 = T2170;
  assign T2170 = 1'h1;
  assign T5859 = T5860 ? 7'h7f : 7'h0;
  assign T5860 = T2167[4'h9];
  assign T2171 = T2093 & T5861;
  assign T5861 = {T5862, T2172};
  assign T2172 = ~ T2168;
  assign T5862 = T5863 ? 7'h7f : 7'h0;
  assign T5863 = T2172[4'h9];
  assign T2173 = T2110 & T2174;
  assign T2174 = 4'h7 == T2109;
  assign T2175 = T2180 | T5864;
  assign T5864 = {T5866, T2176};
  assign T2176 = T5865 & T2177;
  assign T2177 = 9'h80;
  assign T5865 = T2178 ? 9'h1ff : 9'h0;
  assign T2178 = T2179;
  assign T2179 = 1'h1;
  assign T5866 = T5867 ? 8'hff : 8'h0;
  assign T5867 = T2176[4'h8];
  assign T2180 = T2092 & T5868;
  assign T5868 = {T5869, T2181};
  assign T2181 = ~ T2177;
  assign T5869 = T5870 ? 8'hff : 8'h0;
  assign T5870 = T2181[4'h8];
  assign T2182 = T2110 & T2183;
  assign T2183 = 4'h8 == T2109;
  assign T2184 = T2189 | T5871;
  assign T5871 = {T5873, T2185};
  assign T2185 = T5872 & T2186;
  assign T2186 = 8'h40;
  assign T5872 = T2187 ? 8'hff : 8'h0;
  assign T2187 = T2188;
  assign T2188 = 1'h1;
  assign T5873 = T5874 ? 9'h1ff : 9'h0;
  assign T5874 = T2185[3'h7];
  assign T2189 = T2091 & T5875;
  assign T5875 = {T5876, T2190};
  assign T2190 = ~ T2186;
  assign T5876 = T5877 ? 9'h1ff : 9'h0;
  assign T5877 = T2190[3'h7];
  assign T2191 = T2110 & T2192;
  assign T2192 = 4'h9 == T2109;
  assign T2193 = T2198 | T5878;
  assign T5878 = {T5880, T2194};
  assign T2194 = T5879 & T2195;
  assign T2195 = 7'h20;
  assign T5879 = T2196 ? 7'h7f : 7'h0;
  assign T2196 = T2197;
  assign T2197 = 1'h1;
  assign T5880 = T5881 ? 10'h3ff : 10'h0;
  assign T5881 = T2194[3'h6];
  assign T2198 = T2090 & T5882;
  assign T5882 = {T5883, T2199};
  assign T2199 = ~ T2195;
  assign T5883 = T5884 ? 10'h3ff : 10'h0;
  assign T5884 = T2199[3'h6];
  assign T2200 = T2110 & T2201;
  assign T2201 = 4'ha == T2109;
  assign T2202 = T2207 | T5885;
  assign T5885 = {T5887, T2203};
  assign T2203 = T5886 & T2204;
  assign T2204 = 6'h10;
  assign T5886 = T2205 ? 6'h3f : 6'h0;
  assign T2205 = T2206;
  assign T2206 = 1'h1;
  assign T5887 = T5888 ? 11'h7ff : 11'h0;
  assign T5888 = T2203[3'h5];
  assign T2207 = T2089 & T5889;
  assign T5889 = {T5890, T2208};
  assign T2208 = ~ T2204;
  assign T5890 = T5891 ? 11'h7ff : 11'h0;
  assign T5891 = T2208[3'h5];
  assign T2209 = T2110 & T2210;
  assign T2210 = 4'hb == T2109;
  assign T2211 = T2216 | T5892;
  assign T5892 = {T5894, T2212};
  assign T2212 = T5893 & T2213;
  assign T2213 = 5'h8;
  assign T5893 = T2214 ? 5'h1f : 5'h0;
  assign T2214 = T2215;
  assign T2215 = 1'h1;
  assign T5894 = T5895 ? 12'hfff : 12'h0;
  assign T5895 = T2212[3'h4];
  assign T2216 = T2088 & T5896;
  assign T5896 = {T5897, T2217};
  assign T2217 = ~ T2213;
  assign T5897 = T5898 ? 12'hfff : 12'h0;
  assign T5898 = T2217[3'h4];
  assign T2218 = T2110 & T2219;
  assign T2219 = 4'hc == T2109;
  assign T2220 = T2225 | T5899;
  assign T5899 = {T5901, T2221};
  assign T2221 = T5900 & T2222;
  assign T2222 = 4'h4;
  assign T5900 = T2223 ? 4'hf : 4'h0;
  assign T2223 = T2224;
  assign T2224 = 1'h1;
  assign T5901 = T5902 ? 13'h1fff : 13'h0;
  assign T5902 = T2221[2'h3];
  assign T2225 = T2087 & T5903;
  assign T5903 = {T5904, T2226};
  assign T2226 = ~ T2222;
  assign T5904 = T5905 ? 13'h1fff : 13'h0;
  assign T5905 = T2226[2'h3];
  assign T2227 = T2110 & T2228;
  assign T2228 = 4'hd == T2109;
  assign T2229 = T2234 | T5906;
  assign T5906 = {T5908, T2230};
  assign T2230 = T5907 & T2231;
  assign T2231 = 3'h2;
  assign T5907 = T2232 ? 3'h7 : 3'h0;
  assign T2232 = T2233;
  assign T2233 = 1'h1;
  assign T5908 = T5909 ? 14'h3fff : 14'h0;
  assign T5909 = T2230[2'h2];
  assign T2234 = T2086 & T5910;
  assign T5910 = {T5911, T2235};
  assign T2235 = ~ T2231;
  assign T5911 = T5912 ? 14'h3fff : 14'h0;
  assign T5912 = T2235[2'h2];
  assign T2236 = T2110 & T2237;
  assign T2237 = 4'he == T2109;
  assign T2238 = T2243 | T5913;
  assign T5913 = {T5915, T2239};
  assign T2239 = T5914 & T2240;
  assign T2240 = 2'h1;
  assign T5914 = T2241 ? 2'h3 : 2'h0;
  assign T2241 = T2242;
  assign T2242 = 1'h1;
  assign T5915 = T5916 ? 15'h7fff : 15'h0;
  assign T5916 = T2239[1'h1];
  assign T2243 = T2085 & T5917;
  assign T5917 = {T5918, T2244};
  assign T2244 = ~ T2240;
  assign T5918 = T5919 ? 15'h7fff : 15'h0;
  assign T5919 = T2244[1'h1];
  assign T2245 = T2110 & T2246;
  assign T2246 = 4'hf == T2109;
  assign io_V_wire_en_6 = V_wire_en_6;
  assign V_wire_en_6 = T5920;
  assign T5920 = T2247[4'hf:1'h0];
  assign T2247 = T2408 ? T2401 : T2248;
  assign T2248 = T2399 ? T2392 : T2249;
  assign T2249 = T2390 ? T2383 : T2250;
  assign T2250 = T2381 ? T2374 : T2251;
  assign T2251 = T2372 ? T2365 : T2252;
  assign T2252 = T2363 ? T2356 : T2253;
  assign T2253 = T2354 ? T2347 : T2254;
  assign T2254 = T2345 ? T2338 : T2255;
  assign T2255 = T2336 ? T2329 : T2256;
  assign T2256 = T2327 ? T2320 : T2257;
  assign T2257 = T2318 ? T2311 : T2258;
  assign T2258 = T2309 ? T2302 : T2259;
  assign T2259 = T2300 ? T2293 : T2260;
  assign T2260 = T2291 ? T2284 : T2261;
  assign T2261 = T2282 ? T2275 : T2262;
  assign T2262 = T2270 ? T2263 : 17'h0;
  assign T2263 = T2268 | T2264;
  assign T2264 = T5921 & T2265;
  assign T2265 = 17'h8000;
  assign T5921 = T2266 ? 17'h1ffff : 17'h0;
  assign T2266 = T2267;
  assign T2267 = 1'h1;
  assign T2268 = 17'h0 & T2269;
  assign T2269 = ~ T2265;
  assign T2270 = T2273 & T2271;
  assign T2271 = 4'h0 == T2272;
  assign T2272 = LogicBlockModule_6_io_config_V_out[2'h3:1'h0];
  assign T2273 = T2274;
  assign T2274 = LogicBlockModule_6_io_config_V_out[3'h4];
  assign T2275 = T2280 | T5922;
  assign T5922 = {T5924, T2276};
  assign T2276 = T5923 & T2277;
  assign T2277 = 16'h4000;
  assign T5923 = T2278 ? 16'hffff : 16'h0;
  assign T2278 = T2279;
  assign T2279 = 1'h1;
  assign T5924 = T2276[4'hf];
  assign T2280 = T2262 & T5925;
  assign T5925 = {T5926, T2281};
  assign T2281 = ~ T2277;
  assign T5926 = T2281[4'hf];
  assign T2282 = T2273 & T2283;
  assign T2283 = 4'h1 == T2272;
  assign T2284 = T2289 | T5927;
  assign T5927 = {T5929, T2285};
  assign T2285 = T5928 & T2286;
  assign T2286 = 15'h2000;
  assign T5928 = T2287 ? 15'h7fff : 15'h0;
  assign T2287 = T2288;
  assign T2288 = 1'h1;
  assign T5929 = T5930 ? 2'h3 : 2'h0;
  assign T5930 = T2285[4'he];
  assign T2289 = T2261 & T5931;
  assign T5931 = {T5932, T2290};
  assign T2290 = ~ T2286;
  assign T5932 = T5933 ? 2'h3 : 2'h0;
  assign T5933 = T2290[4'he];
  assign T2291 = T2273 & T2292;
  assign T2292 = 4'h2 == T2272;
  assign T2293 = T2298 | T5934;
  assign T5934 = {T5936, T2294};
  assign T2294 = T5935 & T2295;
  assign T2295 = 14'h1000;
  assign T5935 = T2296 ? 14'h3fff : 14'h0;
  assign T2296 = T2297;
  assign T2297 = 1'h1;
  assign T5936 = T5937 ? 3'h7 : 3'h0;
  assign T5937 = T2294[4'hd];
  assign T2298 = T2260 & T5938;
  assign T5938 = {T5939, T2299};
  assign T2299 = ~ T2295;
  assign T5939 = T5940 ? 3'h7 : 3'h0;
  assign T5940 = T2299[4'hd];
  assign T2300 = T2273 & T2301;
  assign T2301 = 4'h3 == T2272;
  assign T2302 = T2307 | T5941;
  assign T5941 = {T5943, T2303};
  assign T2303 = T5942 & T2304;
  assign T2304 = 13'h800;
  assign T5942 = T2305 ? 13'h1fff : 13'h0;
  assign T2305 = T2306;
  assign T2306 = 1'h1;
  assign T5943 = T5944 ? 4'hf : 4'h0;
  assign T5944 = T2303[4'hc];
  assign T2307 = T2259 & T5945;
  assign T5945 = {T5946, T2308};
  assign T2308 = ~ T2304;
  assign T5946 = T5947 ? 4'hf : 4'h0;
  assign T5947 = T2308[4'hc];
  assign T2309 = T2273 & T2310;
  assign T2310 = 4'h4 == T2272;
  assign T2311 = T2316 | T5948;
  assign T5948 = {T5950, T2312};
  assign T2312 = T5949 & T2313;
  assign T2313 = 12'h400;
  assign T5949 = T2314 ? 12'hfff : 12'h0;
  assign T2314 = T2315;
  assign T2315 = 1'h1;
  assign T5950 = T5951 ? 5'h1f : 5'h0;
  assign T5951 = T2312[4'hb];
  assign T2316 = T2258 & T5952;
  assign T5952 = {T5953, T2317};
  assign T2317 = ~ T2313;
  assign T5953 = T5954 ? 5'h1f : 5'h0;
  assign T5954 = T2317[4'hb];
  assign T2318 = T2273 & T2319;
  assign T2319 = 4'h5 == T2272;
  assign T2320 = T2325 | T5955;
  assign T5955 = {T5957, T2321};
  assign T2321 = T5956 & T2322;
  assign T2322 = 11'h200;
  assign T5956 = T2323 ? 11'h7ff : 11'h0;
  assign T2323 = T2324;
  assign T2324 = 1'h1;
  assign T5957 = T5958 ? 6'h3f : 6'h0;
  assign T5958 = T2321[4'ha];
  assign T2325 = T2257 & T5959;
  assign T5959 = {T5960, T2326};
  assign T2326 = ~ T2322;
  assign T5960 = T5961 ? 6'h3f : 6'h0;
  assign T5961 = T2326[4'ha];
  assign T2327 = T2273 & T2328;
  assign T2328 = 4'h6 == T2272;
  assign T2329 = T2334 | T5962;
  assign T5962 = {T5964, T2330};
  assign T2330 = T5963 & T2331;
  assign T2331 = 10'h100;
  assign T5963 = T2332 ? 10'h3ff : 10'h0;
  assign T2332 = T2333;
  assign T2333 = 1'h1;
  assign T5964 = T5965 ? 7'h7f : 7'h0;
  assign T5965 = T2330[4'h9];
  assign T2334 = T2256 & T5966;
  assign T5966 = {T5967, T2335};
  assign T2335 = ~ T2331;
  assign T5967 = T5968 ? 7'h7f : 7'h0;
  assign T5968 = T2335[4'h9];
  assign T2336 = T2273 & T2337;
  assign T2337 = 4'h7 == T2272;
  assign T2338 = T2343 | T5969;
  assign T5969 = {T5971, T2339};
  assign T2339 = T5970 & T2340;
  assign T2340 = 9'h80;
  assign T5970 = T2341 ? 9'h1ff : 9'h0;
  assign T2341 = T2342;
  assign T2342 = 1'h1;
  assign T5971 = T5972 ? 8'hff : 8'h0;
  assign T5972 = T2339[4'h8];
  assign T2343 = T2255 & T5973;
  assign T5973 = {T5974, T2344};
  assign T2344 = ~ T2340;
  assign T5974 = T5975 ? 8'hff : 8'h0;
  assign T5975 = T2344[4'h8];
  assign T2345 = T2273 & T2346;
  assign T2346 = 4'h8 == T2272;
  assign T2347 = T2352 | T5976;
  assign T5976 = {T5978, T2348};
  assign T2348 = T5977 & T2349;
  assign T2349 = 8'h40;
  assign T5977 = T2350 ? 8'hff : 8'h0;
  assign T2350 = T2351;
  assign T2351 = 1'h1;
  assign T5978 = T5979 ? 9'h1ff : 9'h0;
  assign T5979 = T2348[3'h7];
  assign T2352 = T2254 & T5980;
  assign T5980 = {T5981, T2353};
  assign T2353 = ~ T2349;
  assign T5981 = T5982 ? 9'h1ff : 9'h0;
  assign T5982 = T2353[3'h7];
  assign T2354 = T2273 & T2355;
  assign T2355 = 4'h9 == T2272;
  assign T2356 = T2361 | T5983;
  assign T5983 = {T5985, T2357};
  assign T2357 = T5984 & T2358;
  assign T2358 = 7'h20;
  assign T5984 = T2359 ? 7'h7f : 7'h0;
  assign T2359 = T2360;
  assign T2360 = 1'h1;
  assign T5985 = T5986 ? 10'h3ff : 10'h0;
  assign T5986 = T2357[3'h6];
  assign T2361 = T2253 & T5987;
  assign T5987 = {T5988, T2362};
  assign T2362 = ~ T2358;
  assign T5988 = T5989 ? 10'h3ff : 10'h0;
  assign T5989 = T2362[3'h6];
  assign T2363 = T2273 & T2364;
  assign T2364 = 4'ha == T2272;
  assign T2365 = T2370 | T5990;
  assign T5990 = {T5992, T2366};
  assign T2366 = T5991 & T2367;
  assign T2367 = 6'h10;
  assign T5991 = T2368 ? 6'h3f : 6'h0;
  assign T2368 = T2369;
  assign T2369 = 1'h1;
  assign T5992 = T5993 ? 11'h7ff : 11'h0;
  assign T5993 = T2366[3'h5];
  assign T2370 = T2252 & T5994;
  assign T5994 = {T5995, T2371};
  assign T2371 = ~ T2367;
  assign T5995 = T5996 ? 11'h7ff : 11'h0;
  assign T5996 = T2371[3'h5];
  assign T2372 = T2273 & T2373;
  assign T2373 = 4'hb == T2272;
  assign T2374 = T2379 | T5997;
  assign T5997 = {T5999, T2375};
  assign T2375 = T5998 & T2376;
  assign T2376 = 5'h8;
  assign T5998 = T2377 ? 5'h1f : 5'h0;
  assign T2377 = T2378;
  assign T2378 = 1'h1;
  assign T5999 = T6000 ? 12'hfff : 12'h0;
  assign T6000 = T2375[3'h4];
  assign T2379 = T2251 & T6001;
  assign T6001 = {T6002, T2380};
  assign T2380 = ~ T2376;
  assign T6002 = T6003 ? 12'hfff : 12'h0;
  assign T6003 = T2380[3'h4];
  assign T2381 = T2273 & T2382;
  assign T2382 = 4'hc == T2272;
  assign T2383 = T2388 | T6004;
  assign T6004 = {T6006, T2384};
  assign T2384 = T6005 & T2385;
  assign T2385 = 4'h4;
  assign T6005 = T2386 ? 4'hf : 4'h0;
  assign T2386 = T2387;
  assign T2387 = 1'h1;
  assign T6006 = T6007 ? 13'h1fff : 13'h0;
  assign T6007 = T2384[2'h3];
  assign T2388 = T2250 & T6008;
  assign T6008 = {T6009, T2389};
  assign T2389 = ~ T2385;
  assign T6009 = T6010 ? 13'h1fff : 13'h0;
  assign T6010 = T2389[2'h3];
  assign T2390 = T2273 & T2391;
  assign T2391 = 4'hd == T2272;
  assign T2392 = T2397 | T6011;
  assign T6011 = {T6013, T2393};
  assign T2393 = T6012 & T2394;
  assign T2394 = 3'h2;
  assign T6012 = T2395 ? 3'h7 : 3'h0;
  assign T2395 = T2396;
  assign T2396 = 1'h1;
  assign T6013 = T6014 ? 14'h3fff : 14'h0;
  assign T6014 = T2393[2'h2];
  assign T2397 = T2249 & T6015;
  assign T6015 = {T6016, T2398};
  assign T2398 = ~ T2394;
  assign T6016 = T6017 ? 14'h3fff : 14'h0;
  assign T6017 = T2398[2'h2];
  assign T2399 = T2273 & T2400;
  assign T2400 = 4'he == T2272;
  assign T2401 = T2406 | T6018;
  assign T6018 = {T6020, T2402};
  assign T2402 = T6019 & T2403;
  assign T2403 = 2'h1;
  assign T6019 = T2404 ? 2'h3 : 2'h0;
  assign T2404 = T2405;
  assign T2405 = 1'h1;
  assign T6020 = T6021 ? 15'h7fff : 15'h0;
  assign T6021 = T2402[1'h1];
  assign T2406 = T2248 & T6022;
  assign T6022 = {T6023, T2407};
  assign T2407 = ~ T2403;
  assign T6023 = T6024 ? 15'h7fff : 15'h0;
  assign T6024 = T2407[1'h1];
  assign T2408 = T2273 & T2409;
  assign T2409 = 4'hf == T2272;
  assign io_V_wire_en_7 = V_wire_en_7;
  assign V_wire_en_7 = T6025;
  assign T6025 = T2410[4'hf:1'h0];
  assign T2410 = T2571 ? T2564 : T2411;
  assign T2411 = T2562 ? T2555 : T2412;
  assign T2412 = T2553 ? T2546 : T2413;
  assign T2413 = T2544 ? T2537 : T2414;
  assign T2414 = T2535 ? T2528 : T2415;
  assign T2415 = T2526 ? T2519 : T2416;
  assign T2416 = T2517 ? T2510 : T2417;
  assign T2417 = T2508 ? T2501 : T2418;
  assign T2418 = T2499 ? T2492 : T2419;
  assign T2419 = T2490 ? T2483 : T2420;
  assign T2420 = T2481 ? T2474 : T2421;
  assign T2421 = T2472 ? T2465 : T2422;
  assign T2422 = T2463 ? T2456 : T2423;
  assign T2423 = T2454 ? T2447 : T2424;
  assign T2424 = T2445 ? T2438 : T2425;
  assign T2425 = T2433 ? T2426 : 17'h0;
  assign T2426 = T2431 | T2427;
  assign T2427 = T6026 & T2428;
  assign T2428 = 17'h8000;
  assign T6026 = T2429 ? 17'h1ffff : 17'h0;
  assign T2429 = T2430;
  assign T2430 = 1'h1;
  assign T2431 = 17'h0 & T2432;
  assign T2432 = ~ T2428;
  assign T2433 = T2436 & T2434;
  assign T2434 = 4'h0 == T2435;
  assign T2435 = LogicBlockModule_7_io_config_V_out[2'h3:1'h0];
  assign T2436 = T2437;
  assign T2437 = LogicBlockModule_7_io_config_V_out[3'h4];
  assign T2438 = T2443 | T6027;
  assign T6027 = {T6029, T2439};
  assign T2439 = T6028 & T2440;
  assign T2440 = 16'h4000;
  assign T6028 = T2441 ? 16'hffff : 16'h0;
  assign T2441 = T2442;
  assign T2442 = 1'h1;
  assign T6029 = T2439[4'hf];
  assign T2443 = T2425 & T6030;
  assign T6030 = {T6031, T2444};
  assign T2444 = ~ T2440;
  assign T6031 = T2444[4'hf];
  assign T2445 = T2436 & T2446;
  assign T2446 = 4'h1 == T2435;
  assign T2447 = T2452 | T6032;
  assign T6032 = {T6034, T2448};
  assign T2448 = T6033 & T2449;
  assign T2449 = 15'h2000;
  assign T6033 = T2450 ? 15'h7fff : 15'h0;
  assign T2450 = T2451;
  assign T2451 = 1'h1;
  assign T6034 = T6035 ? 2'h3 : 2'h0;
  assign T6035 = T2448[4'he];
  assign T2452 = T2424 & T6036;
  assign T6036 = {T6037, T2453};
  assign T2453 = ~ T2449;
  assign T6037 = T6038 ? 2'h3 : 2'h0;
  assign T6038 = T2453[4'he];
  assign T2454 = T2436 & T2455;
  assign T2455 = 4'h2 == T2435;
  assign T2456 = T2461 | T6039;
  assign T6039 = {T6041, T2457};
  assign T2457 = T6040 & T2458;
  assign T2458 = 14'h1000;
  assign T6040 = T2459 ? 14'h3fff : 14'h0;
  assign T2459 = T2460;
  assign T2460 = 1'h1;
  assign T6041 = T6042 ? 3'h7 : 3'h0;
  assign T6042 = T2457[4'hd];
  assign T2461 = T2423 & T6043;
  assign T6043 = {T6044, T2462};
  assign T2462 = ~ T2458;
  assign T6044 = T6045 ? 3'h7 : 3'h0;
  assign T6045 = T2462[4'hd];
  assign T2463 = T2436 & T2464;
  assign T2464 = 4'h3 == T2435;
  assign T2465 = T2470 | T6046;
  assign T6046 = {T6048, T2466};
  assign T2466 = T6047 & T2467;
  assign T2467 = 13'h800;
  assign T6047 = T2468 ? 13'h1fff : 13'h0;
  assign T2468 = T2469;
  assign T2469 = 1'h1;
  assign T6048 = T6049 ? 4'hf : 4'h0;
  assign T6049 = T2466[4'hc];
  assign T2470 = T2422 & T6050;
  assign T6050 = {T6051, T2471};
  assign T2471 = ~ T2467;
  assign T6051 = T6052 ? 4'hf : 4'h0;
  assign T6052 = T2471[4'hc];
  assign T2472 = T2436 & T2473;
  assign T2473 = 4'h4 == T2435;
  assign T2474 = T2479 | T6053;
  assign T6053 = {T6055, T2475};
  assign T2475 = T6054 & T2476;
  assign T2476 = 12'h400;
  assign T6054 = T2477 ? 12'hfff : 12'h0;
  assign T2477 = T2478;
  assign T2478 = 1'h1;
  assign T6055 = T6056 ? 5'h1f : 5'h0;
  assign T6056 = T2475[4'hb];
  assign T2479 = T2421 & T6057;
  assign T6057 = {T6058, T2480};
  assign T2480 = ~ T2476;
  assign T6058 = T6059 ? 5'h1f : 5'h0;
  assign T6059 = T2480[4'hb];
  assign T2481 = T2436 & T2482;
  assign T2482 = 4'h5 == T2435;
  assign T2483 = T2488 | T6060;
  assign T6060 = {T6062, T2484};
  assign T2484 = T6061 & T2485;
  assign T2485 = 11'h200;
  assign T6061 = T2486 ? 11'h7ff : 11'h0;
  assign T2486 = T2487;
  assign T2487 = 1'h1;
  assign T6062 = T6063 ? 6'h3f : 6'h0;
  assign T6063 = T2484[4'ha];
  assign T2488 = T2420 & T6064;
  assign T6064 = {T6065, T2489};
  assign T2489 = ~ T2485;
  assign T6065 = T6066 ? 6'h3f : 6'h0;
  assign T6066 = T2489[4'ha];
  assign T2490 = T2436 & T2491;
  assign T2491 = 4'h6 == T2435;
  assign T2492 = T2497 | T6067;
  assign T6067 = {T6069, T2493};
  assign T2493 = T6068 & T2494;
  assign T2494 = 10'h100;
  assign T6068 = T2495 ? 10'h3ff : 10'h0;
  assign T2495 = T2496;
  assign T2496 = 1'h1;
  assign T6069 = T6070 ? 7'h7f : 7'h0;
  assign T6070 = T2493[4'h9];
  assign T2497 = T2419 & T6071;
  assign T6071 = {T6072, T2498};
  assign T2498 = ~ T2494;
  assign T6072 = T6073 ? 7'h7f : 7'h0;
  assign T6073 = T2498[4'h9];
  assign T2499 = T2436 & T2500;
  assign T2500 = 4'h7 == T2435;
  assign T2501 = T2506 | T6074;
  assign T6074 = {T6076, T2502};
  assign T2502 = T6075 & T2503;
  assign T2503 = 9'h80;
  assign T6075 = T2504 ? 9'h1ff : 9'h0;
  assign T2504 = T2505;
  assign T2505 = 1'h1;
  assign T6076 = T6077 ? 8'hff : 8'h0;
  assign T6077 = T2502[4'h8];
  assign T2506 = T2418 & T6078;
  assign T6078 = {T6079, T2507};
  assign T2507 = ~ T2503;
  assign T6079 = T6080 ? 8'hff : 8'h0;
  assign T6080 = T2507[4'h8];
  assign T2508 = T2436 & T2509;
  assign T2509 = 4'h8 == T2435;
  assign T2510 = T2515 | T6081;
  assign T6081 = {T6083, T2511};
  assign T2511 = T6082 & T2512;
  assign T2512 = 8'h40;
  assign T6082 = T2513 ? 8'hff : 8'h0;
  assign T2513 = T2514;
  assign T2514 = 1'h1;
  assign T6083 = T6084 ? 9'h1ff : 9'h0;
  assign T6084 = T2511[3'h7];
  assign T2515 = T2417 & T6085;
  assign T6085 = {T6086, T2516};
  assign T2516 = ~ T2512;
  assign T6086 = T6087 ? 9'h1ff : 9'h0;
  assign T6087 = T2516[3'h7];
  assign T2517 = T2436 & T2518;
  assign T2518 = 4'h9 == T2435;
  assign T2519 = T2524 | T6088;
  assign T6088 = {T6090, T2520};
  assign T2520 = T6089 & T2521;
  assign T2521 = 7'h20;
  assign T6089 = T2522 ? 7'h7f : 7'h0;
  assign T2522 = T2523;
  assign T2523 = 1'h1;
  assign T6090 = T6091 ? 10'h3ff : 10'h0;
  assign T6091 = T2520[3'h6];
  assign T2524 = T2416 & T6092;
  assign T6092 = {T6093, T2525};
  assign T2525 = ~ T2521;
  assign T6093 = T6094 ? 10'h3ff : 10'h0;
  assign T6094 = T2525[3'h6];
  assign T2526 = T2436 & T2527;
  assign T2527 = 4'ha == T2435;
  assign T2528 = T2533 | T6095;
  assign T6095 = {T6097, T2529};
  assign T2529 = T6096 & T2530;
  assign T2530 = 6'h10;
  assign T6096 = T2531 ? 6'h3f : 6'h0;
  assign T2531 = T2532;
  assign T2532 = 1'h1;
  assign T6097 = T6098 ? 11'h7ff : 11'h0;
  assign T6098 = T2529[3'h5];
  assign T2533 = T2415 & T6099;
  assign T6099 = {T6100, T2534};
  assign T2534 = ~ T2530;
  assign T6100 = T6101 ? 11'h7ff : 11'h0;
  assign T6101 = T2534[3'h5];
  assign T2535 = T2436 & T2536;
  assign T2536 = 4'hb == T2435;
  assign T2537 = T2542 | T6102;
  assign T6102 = {T6104, T2538};
  assign T2538 = T6103 & T2539;
  assign T2539 = 5'h8;
  assign T6103 = T2540 ? 5'h1f : 5'h0;
  assign T2540 = T2541;
  assign T2541 = 1'h1;
  assign T6104 = T6105 ? 12'hfff : 12'h0;
  assign T6105 = T2538[3'h4];
  assign T2542 = T2414 & T6106;
  assign T6106 = {T6107, T2543};
  assign T2543 = ~ T2539;
  assign T6107 = T6108 ? 12'hfff : 12'h0;
  assign T6108 = T2543[3'h4];
  assign T2544 = T2436 & T2545;
  assign T2545 = 4'hc == T2435;
  assign T2546 = T2551 | T6109;
  assign T6109 = {T6111, T2547};
  assign T2547 = T6110 & T2548;
  assign T2548 = 4'h4;
  assign T6110 = T2549 ? 4'hf : 4'h0;
  assign T2549 = T2550;
  assign T2550 = 1'h1;
  assign T6111 = T6112 ? 13'h1fff : 13'h0;
  assign T6112 = T2547[2'h3];
  assign T2551 = T2413 & T6113;
  assign T6113 = {T6114, T2552};
  assign T2552 = ~ T2548;
  assign T6114 = T6115 ? 13'h1fff : 13'h0;
  assign T6115 = T2552[2'h3];
  assign T2553 = T2436 & T2554;
  assign T2554 = 4'hd == T2435;
  assign T2555 = T2560 | T6116;
  assign T6116 = {T6118, T2556};
  assign T2556 = T6117 & T2557;
  assign T2557 = 3'h2;
  assign T6117 = T2558 ? 3'h7 : 3'h0;
  assign T2558 = T2559;
  assign T2559 = 1'h1;
  assign T6118 = T6119 ? 14'h3fff : 14'h0;
  assign T6119 = T2556[2'h2];
  assign T2560 = T2412 & T6120;
  assign T6120 = {T6121, T2561};
  assign T2561 = ~ T2557;
  assign T6121 = T6122 ? 14'h3fff : 14'h0;
  assign T6122 = T2561[2'h2];
  assign T2562 = T2436 & T2563;
  assign T2563 = 4'he == T2435;
  assign T2564 = T2569 | T6123;
  assign T6123 = {T6125, T2565};
  assign T2565 = T6124 & T2566;
  assign T2566 = 2'h1;
  assign T6124 = T2567 ? 2'h3 : 2'h0;
  assign T2567 = T2568;
  assign T2568 = 1'h1;
  assign T6125 = T6126 ? 15'h7fff : 15'h0;
  assign T6126 = T2565[1'h1];
  assign T2569 = T2411 & T6127;
  assign T6127 = {T6128, T2570};
  assign T2570 = ~ T2566;
  assign T6128 = T6129 ? 15'h7fff : 15'h0;
  assign T6129 = T2570[1'h1];
  assign T2571 = T2436 & T2572;
  assign T2572 = 4'hf == T2435;
  assign io_V_wire_en_8 = V_wire_en_8;
  assign V_wire_en_8 = T6130;
  assign T6130 = T2573[4'hf:1'h0];
  assign T2573 = T2734 ? T2727 : T2574;
  assign T2574 = T2725 ? T2718 : T2575;
  assign T2575 = T2716 ? T2709 : T2576;
  assign T2576 = T2707 ? T2700 : T2577;
  assign T2577 = T2698 ? T2691 : T2578;
  assign T2578 = T2689 ? T2682 : T2579;
  assign T2579 = T2680 ? T2673 : T2580;
  assign T2580 = T2671 ? T2664 : T2581;
  assign T2581 = T2662 ? T2655 : T2582;
  assign T2582 = T2653 ? T2646 : T2583;
  assign T2583 = T2644 ? T2637 : T2584;
  assign T2584 = T2635 ? T2628 : T2585;
  assign T2585 = T2626 ? T2619 : T2586;
  assign T2586 = T2617 ? T2610 : T2587;
  assign T2587 = T2608 ? T2601 : T2588;
  assign T2588 = T2596 ? T2589 : 17'h0;
  assign T2589 = T2594 | T2590;
  assign T2590 = T6131 & T2591;
  assign T2591 = 17'h8000;
  assign T6131 = T2592 ? 17'h1ffff : 17'h0;
  assign T2592 = T2593;
  assign T2593 = 1'h1;
  assign T2594 = 17'h0 & T2595;
  assign T2595 = ~ T2591;
  assign T2596 = T2599 & T2597;
  assign T2597 = 4'h0 == T2598;
  assign T2598 = LogicBlockModule_8_io_config_V_out[2'h3:1'h0];
  assign T2599 = T2600;
  assign T2600 = LogicBlockModule_8_io_config_V_out[3'h4];
  assign T2601 = T2606 | T6132;
  assign T6132 = {T6134, T2602};
  assign T2602 = T6133 & T2603;
  assign T2603 = 16'h4000;
  assign T6133 = T2604 ? 16'hffff : 16'h0;
  assign T2604 = T2605;
  assign T2605 = 1'h1;
  assign T6134 = T2602[4'hf];
  assign T2606 = T2588 & T6135;
  assign T6135 = {T6136, T2607};
  assign T2607 = ~ T2603;
  assign T6136 = T2607[4'hf];
  assign T2608 = T2599 & T2609;
  assign T2609 = 4'h1 == T2598;
  assign T2610 = T2615 | T6137;
  assign T6137 = {T6139, T2611};
  assign T2611 = T6138 & T2612;
  assign T2612 = 15'h2000;
  assign T6138 = T2613 ? 15'h7fff : 15'h0;
  assign T2613 = T2614;
  assign T2614 = 1'h1;
  assign T6139 = T6140 ? 2'h3 : 2'h0;
  assign T6140 = T2611[4'he];
  assign T2615 = T2587 & T6141;
  assign T6141 = {T6142, T2616};
  assign T2616 = ~ T2612;
  assign T6142 = T6143 ? 2'h3 : 2'h0;
  assign T6143 = T2616[4'he];
  assign T2617 = T2599 & T2618;
  assign T2618 = 4'h2 == T2598;
  assign T2619 = T2624 | T6144;
  assign T6144 = {T6146, T2620};
  assign T2620 = T6145 & T2621;
  assign T2621 = 14'h1000;
  assign T6145 = T2622 ? 14'h3fff : 14'h0;
  assign T2622 = T2623;
  assign T2623 = 1'h1;
  assign T6146 = T6147 ? 3'h7 : 3'h0;
  assign T6147 = T2620[4'hd];
  assign T2624 = T2586 & T6148;
  assign T6148 = {T6149, T2625};
  assign T2625 = ~ T2621;
  assign T6149 = T6150 ? 3'h7 : 3'h0;
  assign T6150 = T2625[4'hd];
  assign T2626 = T2599 & T2627;
  assign T2627 = 4'h3 == T2598;
  assign T2628 = T2633 | T6151;
  assign T6151 = {T6153, T2629};
  assign T2629 = T6152 & T2630;
  assign T2630 = 13'h800;
  assign T6152 = T2631 ? 13'h1fff : 13'h0;
  assign T2631 = T2632;
  assign T2632 = 1'h1;
  assign T6153 = T6154 ? 4'hf : 4'h0;
  assign T6154 = T2629[4'hc];
  assign T2633 = T2585 & T6155;
  assign T6155 = {T6156, T2634};
  assign T2634 = ~ T2630;
  assign T6156 = T6157 ? 4'hf : 4'h0;
  assign T6157 = T2634[4'hc];
  assign T2635 = T2599 & T2636;
  assign T2636 = 4'h4 == T2598;
  assign T2637 = T2642 | T6158;
  assign T6158 = {T6160, T2638};
  assign T2638 = T6159 & T2639;
  assign T2639 = 12'h400;
  assign T6159 = T2640 ? 12'hfff : 12'h0;
  assign T2640 = T2641;
  assign T2641 = 1'h1;
  assign T6160 = T6161 ? 5'h1f : 5'h0;
  assign T6161 = T2638[4'hb];
  assign T2642 = T2584 & T6162;
  assign T6162 = {T6163, T2643};
  assign T2643 = ~ T2639;
  assign T6163 = T6164 ? 5'h1f : 5'h0;
  assign T6164 = T2643[4'hb];
  assign T2644 = T2599 & T2645;
  assign T2645 = 4'h5 == T2598;
  assign T2646 = T2651 | T6165;
  assign T6165 = {T6167, T2647};
  assign T2647 = T6166 & T2648;
  assign T2648 = 11'h200;
  assign T6166 = T2649 ? 11'h7ff : 11'h0;
  assign T2649 = T2650;
  assign T2650 = 1'h1;
  assign T6167 = T6168 ? 6'h3f : 6'h0;
  assign T6168 = T2647[4'ha];
  assign T2651 = T2583 & T6169;
  assign T6169 = {T6170, T2652};
  assign T2652 = ~ T2648;
  assign T6170 = T6171 ? 6'h3f : 6'h0;
  assign T6171 = T2652[4'ha];
  assign T2653 = T2599 & T2654;
  assign T2654 = 4'h6 == T2598;
  assign T2655 = T2660 | T6172;
  assign T6172 = {T6174, T2656};
  assign T2656 = T6173 & T2657;
  assign T2657 = 10'h100;
  assign T6173 = T2658 ? 10'h3ff : 10'h0;
  assign T2658 = T2659;
  assign T2659 = 1'h1;
  assign T6174 = T6175 ? 7'h7f : 7'h0;
  assign T6175 = T2656[4'h9];
  assign T2660 = T2582 & T6176;
  assign T6176 = {T6177, T2661};
  assign T2661 = ~ T2657;
  assign T6177 = T6178 ? 7'h7f : 7'h0;
  assign T6178 = T2661[4'h9];
  assign T2662 = T2599 & T2663;
  assign T2663 = 4'h7 == T2598;
  assign T2664 = T2669 | T6179;
  assign T6179 = {T6181, T2665};
  assign T2665 = T6180 & T2666;
  assign T2666 = 9'h80;
  assign T6180 = T2667 ? 9'h1ff : 9'h0;
  assign T2667 = T2668;
  assign T2668 = 1'h1;
  assign T6181 = T6182 ? 8'hff : 8'h0;
  assign T6182 = T2665[4'h8];
  assign T2669 = T2581 & T6183;
  assign T6183 = {T6184, T2670};
  assign T2670 = ~ T2666;
  assign T6184 = T6185 ? 8'hff : 8'h0;
  assign T6185 = T2670[4'h8];
  assign T2671 = T2599 & T2672;
  assign T2672 = 4'h8 == T2598;
  assign T2673 = T2678 | T6186;
  assign T6186 = {T6188, T2674};
  assign T2674 = T6187 & T2675;
  assign T2675 = 8'h40;
  assign T6187 = T2676 ? 8'hff : 8'h0;
  assign T2676 = T2677;
  assign T2677 = 1'h1;
  assign T6188 = T6189 ? 9'h1ff : 9'h0;
  assign T6189 = T2674[3'h7];
  assign T2678 = T2580 & T6190;
  assign T6190 = {T6191, T2679};
  assign T2679 = ~ T2675;
  assign T6191 = T6192 ? 9'h1ff : 9'h0;
  assign T6192 = T2679[3'h7];
  assign T2680 = T2599 & T2681;
  assign T2681 = 4'h9 == T2598;
  assign T2682 = T2687 | T6193;
  assign T6193 = {T6195, T2683};
  assign T2683 = T6194 & T2684;
  assign T2684 = 7'h20;
  assign T6194 = T2685 ? 7'h7f : 7'h0;
  assign T2685 = T2686;
  assign T2686 = 1'h1;
  assign T6195 = T6196 ? 10'h3ff : 10'h0;
  assign T6196 = T2683[3'h6];
  assign T2687 = T2579 & T6197;
  assign T6197 = {T6198, T2688};
  assign T2688 = ~ T2684;
  assign T6198 = T6199 ? 10'h3ff : 10'h0;
  assign T6199 = T2688[3'h6];
  assign T2689 = T2599 & T2690;
  assign T2690 = 4'ha == T2598;
  assign T2691 = T2696 | T6200;
  assign T6200 = {T6202, T2692};
  assign T2692 = T6201 & T2693;
  assign T2693 = 6'h10;
  assign T6201 = T2694 ? 6'h3f : 6'h0;
  assign T2694 = T2695;
  assign T2695 = 1'h1;
  assign T6202 = T6203 ? 11'h7ff : 11'h0;
  assign T6203 = T2692[3'h5];
  assign T2696 = T2578 & T6204;
  assign T6204 = {T6205, T2697};
  assign T2697 = ~ T2693;
  assign T6205 = T6206 ? 11'h7ff : 11'h0;
  assign T6206 = T2697[3'h5];
  assign T2698 = T2599 & T2699;
  assign T2699 = 4'hb == T2598;
  assign T2700 = T2705 | T6207;
  assign T6207 = {T6209, T2701};
  assign T2701 = T6208 & T2702;
  assign T2702 = 5'h8;
  assign T6208 = T2703 ? 5'h1f : 5'h0;
  assign T2703 = T2704;
  assign T2704 = 1'h1;
  assign T6209 = T6210 ? 12'hfff : 12'h0;
  assign T6210 = T2701[3'h4];
  assign T2705 = T2577 & T6211;
  assign T6211 = {T6212, T2706};
  assign T2706 = ~ T2702;
  assign T6212 = T6213 ? 12'hfff : 12'h0;
  assign T6213 = T2706[3'h4];
  assign T2707 = T2599 & T2708;
  assign T2708 = 4'hc == T2598;
  assign T2709 = T2714 | T6214;
  assign T6214 = {T6216, T2710};
  assign T2710 = T6215 & T2711;
  assign T2711 = 4'h4;
  assign T6215 = T2712 ? 4'hf : 4'h0;
  assign T2712 = T2713;
  assign T2713 = 1'h1;
  assign T6216 = T6217 ? 13'h1fff : 13'h0;
  assign T6217 = T2710[2'h3];
  assign T2714 = T2576 & T6218;
  assign T6218 = {T6219, T2715};
  assign T2715 = ~ T2711;
  assign T6219 = T6220 ? 13'h1fff : 13'h0;
  assign T6220 = T2715[2'h3];
  assign T2716 = T2599 & T2717;
  assign T2717 = 4'hd == T2598;
  assign T2718 = T2723 | T6221;
  assign T6221 = {T6223, T2719};
  assign T2719 = T6222 & T2720;
  assign T2720 = 3'h2;
  assign T6222 = T2721 ? 3'h7 : 3'h0;
  assign T2721 = T2722;
  assign T2722 = 1'h1;
  assign T6223 = T6224 ? 14'h3fff : 14'h0;
  assign T6224 = T2719[2'h2];
  assign T2723 = T2575 & T6225;
  assign T6225 = {T6226, T2724};
  assign T2724 = ~ T2720;
  assign T6226 = T6227 ? 14'h3fff : 14'h0;
  assign T6227 = T2724[2'h2];
  assign T2725 = T2599 & T2726;
  assign T2726 = 4'he == T2598;
  assign T2727 = T2732 | T6228;
  assign T6228 = {T6230, T2728};
  assign T2728 = T6229 & T2729;
  assign T2729 = 2'h1;
  assign T6229 = T2730 ? 2'h3 : 2'h0;
  assign T2730 = T2731;
  assign T2731 = 1'h1;
  assign T6230 = T6231 ? 15'h7fff : 15'h0;
  assign T6231 = T2728[1'h1];
  assign T2732 = T2574 & T6232;
  assign T6232 = {T6233, T2733};
  assign T2733 = ~ T2729;
  assign T6233 = T6234 ? 15'h7fff : 15'h0;
  assign T6234 = T2733[1'h1];
  assign T2734 = T2599 & T2735;
  assign T2735 = 4'hf == T2598;
  assign io_V_wire_en_9 = V_wire_en_9;
  assign V_wire_en_9 = T6235;
  assign T6235 = T2736[4'hf:1'h0];
  assign T2736 = T2897 ? T2890 : T2737;
  assign T2737 = T2888 ? T2881 : T2738;
  assign T2738 = T2879 ? T2872 : T2739;
  assign T2739 = T2870 ? T2863 : T2740;
  assign T2740 = T2861 ? T2854 : T2741;
  assign T2741 = T2852 ? T2845 : T2742;
  assign T2742 = T2843 ? T2836 : T2743;
  assign T2743 = T2834 ? T2827 : T2744;
  assign T2744 = T2825 ? T2818 : T2745;
  assign T2745 = T2816 ? T2809 : T2746;
  assign T2746 = T2807 ? T2800 : T2747;
  assign T2747 = T2798 ? T2791 : T2748;
  assign T2748 = T2789 ? T2782 : T2749;
  assign T2749 = T2780 ? T2773 : T2750;
  assign T2750 = T2771 ? T2764 : T2751;
  assign T2751 = T2759 ? T2752 : 17'h0;
  assign T2752 = T2757 | T2753;
  assign T2753 = T6236 & T2754;
  assign T2754 = 17'h8000;
  assign T6236 = T2755 ? 17'h1ffff : 17'h0;
  assign T2755 = T2756;
  assign T2756 = 1'h1;
  assign T2757 = 17'h0 & T2758;
  assign T2758 = ~ T2754;
  assign T2759 = T2762 & T2760;
  assign T2760 = 4'h0 == T2761;
  assign T2761 = LogicBlockModule_9_io_config_V_out[2'h3:1'h0];
  assign T2762 = T2763;
  assign T2763 = LogicBlockModule_9_io_config_V_out[3'h4];
  assign T2764 = T2769 | T6237;
  assign T6237 = {T6239, T2765};
  assign T2765 = T6238 & T2766;
  assign T2766 = 16'h4000;
  assign T6238 = T2767 ? 16'hffff : 16'h0;
  assign T2767 = T2768;
  assign T2768 = 1'h1;
  assign T6239 = T2765[4'hf];
  assign T2769 = T2751 & T6240;
  assign T6240 = {T6241, T2770};
  assign T2770 = ~ T2766;
  assign T6241 = T2770[4'hf];
  assign T2771 = T2762 & T2772;
  assign T2772 = 4'h1 == T2761;
  assign T2773 = T2778 | T6242;
  assign T6242 = {T6244, T2774};
  assign T2774 = T6243 & T2775;
  assign T2775 = 15'h2000;
  assign T6243 = T2776 ? 15'h7fff : 15'h0;
  assign T2776 = T2777;
  assign T2777 = 1'h1;
  assign T6244 = T6245 ? 2'h3 : 2'h0;
  assign T6245 = T2774[4'he];
  assign T2778 = T2750 & T6246;
  assign T6246 = {T6247, T2779};
  assign T2779 = ~ T2775;
  assign T6247 = T6248 ? 2'h3 : 2'h0;
  assign T6248 = T2779[4'he];
  assign T2780 = T2762 & T2781;
  assign T2781 = 4'h2 == T2761;
  assign T2782 = T2787 | T6249;
  assign T6249 = {T6251, T2783};
  assign T2783 = T6250 & T2784;
  assign T2784 = 14'h1000;
  assign T6250 = T2785 ? 14'h3fff : 14'h0;
  assign T2785 = T2786;
  assign T2786 = 1'h1;
  assign T6251 = T6252 ? 3'h7 : 3'h0;
  assign T6252 = T2783[4'hd];
  assign T2787 = T2749 & T6253;
  assign T6253 = {T6254, T2788};
  assign T2788 = ~ T2784;
  assign T6254 = T6255 ? 3'h7 : 3'h0;
  assign T6255 = T2788[4'hd];
  assign T2789 = T2762 & T2790;
  assign T2790 = 4'h3 == T2761;
  assign T2791 = T2796 | T6256;
  assign T6256 = {T6258, T2792};
  assign T2792 = T6257 & T2793;
  assign T2793 = 13'h800;
  assign T6257 = T2794 ? 13'h1fff : 13'h0;
  assign T2794 = T2795;
  assign T2795 = 1'h1;
  assign T6258 = T6259 ? 4'hf : 4'h0;
  assign T6259 = T2792[4'hc];
  assign T2796 = T2748 & T6260;
  assign T6260 = {T6261, T2797};
  assign T2797 = ~ T2793;
  assign T6261 = T6262 ? 4'hf : 4'h0;
  assign T6262 = T2797[4'hc];
  assign T2798 = T2762 & T2799;
  assign T2799 = 4'h4 == T2761;
  assign T2800 = T2805 | T6263;
  assign T6263 = {T6265, T2801};
  assign T2801 = T6264 & T2802;
  assign T2802 = 12'h400;
  assign T6264 = T2803 ? 12'hfff : 12'h0;
  assign T2803 = T2804;
  assign T2804 = 1'h1;
  assign T6265 = T6266 ? 5'h1f : 5'h0;
  assign T6266 = T2801[4'hb];
  assign T2805 = T2747 & T6267;
  assign T6267 = {T6268, T2806};
  assign T2806 = ~ T2802;
  assign T6268 = T6269 ? 5'h1f : 5'h0;
  assign T6269 = T2806[4'hb];
  assign T2807 = T2762 & T2808;
  assign T2808 = 4'h5 == T2761;
  assign T2809 = T2814 | T6270;
  assign T6270 = {T6272, T2810};
  assign T2810 = T6271 & T2811;
  assign T2811 = 11'h200;
  assign T6271 = T2812 ? 11'h7ff : 11'h0;
  assign T2812 = T2813;
  assign T2813 = 1'h1;
  assign T6272 = T6273 ? 6'h3f : 6'h0;
  assign T6273 = T2810[4'ha];
  assign T2814 = T2746 & T6274;
  assign T6274 = {T6275, T2815};
  assign T2815 = ~ T2811;
  assign T6275 = T6276 ? 6'h3f : 6'h0;
  assign T6276 = T2815[4'ha];
  assign T2816 = T2762 & T2817;
  assign T2817 = 4'h6 == T2761;
  assign T2818 = T2823 | T6277;
  assign T6277 = {T6279, T2819};
  assign T2819 = T6278 & T2820;
  assign T2820 = 10'h100;
  assign T6278 = T2821 ? 10'h3ff : 10'h0;
  assign T2821 = T2822;
  assign T2822 = 1'h1;
  assign T6279 = T6280 ? 7'h7f : 7'h0;
  assign T6280 = T2819[4'h9];
  assign T2823 = T2745 & T6281;
  assign T6281 = {T6282, T2824};
  assign T2824 = ~ T2820;
  assign T6282 = T6283 ? 7'h7f : 7'h0;
  assign T6283 = T2824[4'h9];
  assign T2825 = T2762 & T2826;
  assign T2826 = 4'h7 == T2761;
  assign T2827 = T2832 | T6284;
  assign T6284 = {T6286, T2828};
  assign T2828 = T6285 & T2829;
  assign T2829 = 9'h80;
  assign T6285 = T2830 ? 9'h1ff : 9'h0;
  assign T2830 = T2831;
  assign T2831 = 1'h1;
  assign T6286 = T6287 ? 8'hff : 8'h0;
  assign T6287 = T2828[4'h8];
  assign T2832 = T2744 & T6288;
  assign T6288 = {T6289, T2833};
  assign T2833 = ~ T2829;
  assign T6289 = T6290 ? 8'hff : 8'h0;
  assign T6290 = T2833[4'h8];
  assign T2834 = T2762 & T2835;
  assign T2835 = 4'h8 == T2761;
  assign T2836 = T2841 | T6291;
  assign T6291 = {T6293, T2837};
  assign T2837 = T6292 & T2838;
  assign T2838 = 8'h40;
  assign T6292 = T2839 ? 8'hff : 8'h0;
  assign T2839 = T2840;
  assign T2840 = 1'h1;
  assign T6293 = T6294 ? 9'h1ff : 9'h0;
  assign T6294 = T2837[3'h7];
  assign T2841 = T2743 & T6295;
  assign T6295 = {T6296, T2842};
  assign T2842 = ~ T2838;
  assign T6296 = T6297 ? 9'h1ff : 9'h0;
  assign T6297 = T2842[3'h7];
  assign T2843 = T2762 & T2844;
  assign T2844 = 4'h9 == T2761;
  assign T2845 = T2850 | T6298;
  assign T6298 = {T6300, T2846};
  assign T2846 = T6299 & T2847;
  assign T2847 = 7'h20;
  assign T6299 = T2848 ? 7'h7f : 7'h0;
  assign T2848 = T2849;
  assign T2849 = 1'h1;
  assign T6300 = T6301 ? 10'h3ff : 10'h0;
  assign T6301 = T2846[3'h6];
  assign T2850 = T2742 & T6302;
  assign T6302 = {T6303, T2851};
  assign T2851 = ~ T2847;
  assign T6303 = T6304 ? 10'h3ff : 10'h0;
  assign T6304 = T2851[3'h6];
  assign T2852 = T2762 & T2853;
  assign T2853 = 4'ha == T2761;
  assign T2854 = T2859 | T6305;
  assign T6305 = {T6307, T2855};
  assign T2855 = T6306 & T2856;
  assign T2856 = 6'h10;
  assign T6306 = T2857 ? 6'h3f : 6'h0;
  assign T2857 = T2858;
  assign T2858 = 1'h1;
  assign T6307 = T6308 ? 11'h7ff : 11'h0;
  assign T6308 = T2855[3'h5];
  assign T2859 = T2741 & T6309;
  assign T6309 = {T6310, T2860};
  assign T2860 = ~ T2856;
  assign T6310 = T6311 ? 11'h7ff : 11'h0;
  assign T6311 = T2860[3'h5];
  assign T2861 = T2762 & T2862;
  assign T2862 = 4'hb == T2761;
  assign T2863 = T2868 | T6312;
  assign T6312 = {T6314, T2864};
  assign T2864 = T6313 & T2865;
  assign T2865 = 5'h8;
  assign T6313 = T2866 ? 5'h1f : 5'h0;
  assign T2866 = T2867;
  assign T2867 = 1'h1;
  assign T6314 = T6315 ? 12'hfff : 12'h0;
  assign T6315 = T2864[3'h4];
  assign T2868 = T2740 & T6316;
  assign T6316 = {T6317, T2869};
  assign T2869 = ~ T2865;
  assign T6317 = T6318 ? 12'hfff : 12'h0;
  assign T6318 = T2869[3'h4];
  assign T2870 = T2762 & T2871;
  assign T2871 = 4'hc == T2761;
  assign T2872 = T2877 | T6319;
  assign T6319 = {T6321, T2873};
  assign T2873 = T6320 & T2874;
  assign T2874 = 4'h4;
  assign T6320 = T2875 ? 4'hf : 4'h0;
  assign T2875 = T2876;
  assign T2876 = 1'h1;
  assign T6321 = T6322 ? 13'h1fff : 13'h0;
  assign T6322 = T2873[2'h3];
  assign T2877 = T2739 & T6323;
  assign T6323 = {T6324, T2878};
  assign T2878 = ~ T2874;
  assign T6324 = T6325 ? 13'h1fff : 13'h0;
  assign T6325 = T2878[2'h3];
  assign T2879 = T2762 & T2880;
  assign T2880 = 4'hd == T2761;
  assign T2881 = T2886 | T6326;
  assign T6326 = {T6328, T2882};
  assign T2882 = T6327 & T2883;
  assign T2883 = 3'h2;
  assign T6327 = T2884 ? 3'h7 : 3'h0;
  assign T2884 = T2885;
  assign T2885 = 1'h1;
  assign T6328 = T6329 ? 14'h3fff : 14'h0;
  assign T6329 = T2882[2'h2];
  assign T2886 = T2738 & T6330;
  assign T6330 = {T6331, T2887};
  assign T2887 = ~ T2883;
  assign T6331 = T6332 ? 14'h3fff : 14'h0;
  assign T6332 = T2887[2'h2];
  assign T2888 = T2762 & T2889;
  assign T2889 = 4'he == T2761;
  assign T2890 = T2895 | T6333;
  assign T6333 = {T6335, T2891};
  assign T2891 = T6334 & T2892;
  assign T2892 = 2'h1;
  assign T6334 = T2893 ? 2'h3 : 2'h0;
  assign T2893 = T2894;
  assign T2894 = 1'h1;
  assign T6335 = T6336 ? 15'h7fff : 15'h0;
  assign T6336 = T2891[1'h1];
  assign T2895 = T2737 & T6337;
  assign T6337 = {T6338, T2896};
  assign T2896 = ~ T2892;
  assign T6338 = T6339 ? 15'h7fff : 15'h0;
  assign T6339 = T2896[1'h1];
  assign T2897 = T2762 & T2898;
  assign T2898 = 4'hf == T2761;
  assign io_V_wire_en_10 = V_wire_en_10;
  assign V_wire_en_10 = T6340;
  assign T6340 = T2899[4'hf:1'h0];
  assign T2899 = T3060 ? T3053 : T2900;
  assign T2900 = T3051 ? T3044 : T2901;
  assign T2901 = T3042 ? T3035 : T2902;
  assign T2902 = T3033 ? T3026 : T2903;
  assign T2903 = T3024 ? T3017 : T2904;
  assign T2904 = T3015 ? T3008 : T2905;
  assign T2905 = T3006 ? T2999 : T2906;
  assign T2906 = T2997 ? T2990 : T2907;
  assign T2907 = T2988 ? T2981 : T2908;
  assign T2908 = T2979 ? T2972 : T2909;
  assign T2909 = T2970 ? T2963 : T2910;
  assign T2910 = T2961 ? T2954 : T2911;
  assign T2911 = T2952 ? T2945 : T2912;
  assign T2912 = T2943 ? T2936 : T2913;
  assign T2913 = T2934 ? T2927 : T2914;
  assign T2914 = T2922 ? T2915 : 17'h0;
  assign T2915 = T2920 | T2916;
  assign T2916 = T6341 & T2917;
  assign T2917 = 17'h8000;
  assign T6341 = T2918 ? 17'h1ffff : 17'h0;
  assign T2918 = T2919;
  assign T2919 = 1'h1;
  assign T2920 = 17'h0 & T2921;
  assign T2921 = ~ T2917;
  assign T2922 = T2925 & T2923;
  assign T2923 = 4'h0 == T2924;
  assign T2924 = LogicBlockModule_10_io_config_V_out[2'h3:1'h0];
  assign T2925 = T2926;
  assign T2926 = LogicBlockModule_10_io_config_V_out[3'h4];
  assign T2927 = T2932 | T6342;
  assign T6342 = {T6344, T2928};
  assign T2928 = T6343 & T2929;
  assign T2929 = 16'h4000;
  assign T6343 = T2930 ? 16'hffff : 16'h0;
  assign T2930 = T2931;
  assign T2931 = 1'h1;
  assign T6344 = T2928[4'hf];
  assign T2932 = T2914 & T6345;
  assign T6345 = {T6346, T2933};
  assign T2933 = ~ T2929;
  assign T6346 = T2933[4'hf];
  assign T2934 = T2925 & T2935;
  assign T2935 = 4'h1 == T2924;
  assign T2936 = T2941 | T6347;
  assign T6347 = {T6349, T2937};
  assign T2937 = T6348 & T2938;
  assign T2938 = 15'h2000;
  assign T6348 = T2939 ? 15'h7fff : 15'h0;
  assign T2939 = T2940;
  assign T2940 = 1'h1;
  assign T6349 = T6350 ? 2'h3 : 2'h0;
  assign T6350 = T2937[4'he];
  assign T2941 = T2913 & T6351;
  assign T6351 = {T6352, T2942};
  assign T2942 = ~ T2938;
  assign T6352 = T6353 ? 2'h3 : 2'h0;
  assign T6353 = T2942[4'he];
  assign T2943 = T2925 & T2944;
  assign T2944 = 4'h2 == T2924;
  assign T2945 = T2950 | T6354;
  assign T6354 = {T6356, T2946};
  assign T2946 = T6355 & T2947;
  assign T2947 = 14'h1000;
  assign T6355 = T2948 ? 14'h3fff : 14'h0;
  assign T2948 = T2949;
  assign T2949 = 1'h1;
  assign T6356 = T6357 ? 3'h7 : 3'h0;
  assign T6357 = T2946[4'hd];
  assign T2950 = T2912 & T6358;
  assign T6358 = {T6359, T2951};
  assign T2951 = ~ T2947;
  assign T6359 = T6360 ? 3'h7 : 3'h0;
  assign T6360 = T2951[4'hd];
  assign T2952 = T2925 & T2953;
  assign T2953 = 4'h3 == T2924;
  assign T2954 = T2959 | T6361;
  assign T6361 = {T6363, T2955};
  assign T2955 = T6362 & T2956;
  assign T2956 = 13'h800;
  assign T6362 = T2957 ? 13'h1fff : 13'h0;
  assign T2957 = T2958;
  assign T2958 = 1'h1;
  assign T6363 = T6364 ? 4'hf : 4'h0;
  assign T6364 = T2955[4'hc];
  assign T2959 = T2911 & T6365;
  assign T6365 = {T6366, T2960};
  assign T2960 = ~ T2956;
  assign T6366 = T6367 ? 4'hf : 4'h0;
  assign T6367 = T2960[4'hc];
  assign T2961 = T2925 & T2962;
  assign T2962 = 4'h4 == T2924;
  assign T2963 = T2968 | T6368;
  assign T6368 = {T6370, T2964};
  assign T2964 = T6369 & T2965;
  assign T2965 = 12'h400;
  assign T6369 = T2966 ? 12'hfff : 12'h0;
  assign T2966 = T2967;
  assign T2967 = 1'h1;
  assign T6370 = T6371 ? 5'h1f : 5'h0;
  assign T6371 = T2964[4'hb];
  assign T2968 = T2910 & T6372;
  assign T6372 = {T6373, T2969};
  assign T2969 = ~ T2965;
  assign T6373 = T6374 ? 5'h1f : 5'h0;
  assign T6374 = T2969[4'hb];
  assign T2970 = T2925 & T2971;
  assign T2971 = 4'h5 == T2924;
  assign T2972 = T2977 | T6375;
  assign T6375 = {T6377, T2973};
  assign T2973 = T6376 & T2974;
  assign T2974 = 11'h200;
  assign T6376 = T2975 ? 11'h7ff : 11'h0;
  assign T2975 = T2976;
  assign T2976 = 1'h1;
  assign T6377 = T6378 ? 6'h3f : 6'h0;
  assign T6378 = T2973[4'ha];
  assign T2977 = T2909 & T6379;
  assign T6379 = {T6380, T2978};
  assign T2978 = ~ T2974;
  assign T6380 = T6381 ? 6'h3f : 6'h0;
  assign T6381 = T2978[4'ha];
  assign T2979 = T2925 & T2980;
  assign T2980 = 4'h6 == T2924;
  assign T2981 = T2986 | T6382;
  assign T6382 = {T6384, T2982};
  assign T2982 = T6383 & T2983;
  assign T2983 = 10'h100;
  assign T6383 = T2984 ? 10'h3ff : 10'h0;
  assign T2984 = T2985;
  assign T2985 = 1'h1;
  assign T6384 = T6385 ? 7'h7f : 7'h0;
  assign T6385 = T2982[4'h9];
  assign T2986 = T2908 & T6386;
  assign T6386 = {T6387, T2987};
  assign T2987 = ~ T2983;
  assign T6387 = T6388 ? 7'h7f : 7'h0;
  assign T6388 = T2987[4'h9];
  assign T2988 = T2925 & T2989;
  assign T2989 = 4'h7 == T2924;
  assign T2990 = T2995 | T6389;
  assign T6389 = {T6391, T2991};
  assign T2991 = T6390 & T2992;
  assign T2992 = 9'h80;
  assign T6390 = T2993 ? 9'h1ff : 9'h0;
  assign T2993 = T2994;
  assign T2994 = 1'h1;
  assign T6391 = T6392 ? 8'hff : 8'h0;
  assign T6392 = T2991[4'h8];
  assign T2995 = T2907 & T6393;
  assign T6393 = {T6394, T2996};
  assign T2996 = ~ T2992;
  assign T6394 = T6395 ? 8'hff : 8'h0;
  assign T6395 = T2996[4'h8];
  assign T2997 = T2925 & T2998;
  assign T2998 = 4'h8 == T2924;
  assign T2999 = T3004 | T6396;
  assign T6396 = {T6398, T3000};
  assign T3000 = T6397 & T3001;
  assign T3001 = 8'h40;
  assign T6397 = T3002 ? 8'hff : 8'h0;
  assign T3002 = T3003;
  assign T3003 = 1'h1;
  assign T6398 = T6399 ? 9'h1ff : 9'h0;
  assign T6399 = T3000[3'h7];
  assign T3004 = T2906 & T6400;
  assign T6400 = {T6401, T3005};
  assign T3005 = ~ T3001;
  assign T6401 = T6402 ? 9'h1ff : 9'h0;
  assign T6402 = T3005[3'h7];
  assign T3006 = T2925 & T3007;
  assign T3007 = 4'h9 == T2924;
  assign T3008 = T3013 | T6403;
  assign T6403 = {T6405, T3009};
  assign T3009 = T6404 & T3010;
  assign T3010 = 7'h20;
  assign T6404 = T3011 ? 7'h7f : 7'h0;
  assign T3011 = T3012;
  assign T3012 = 1'h1;
  assign T6405 = T6406 ? 10'h3ff : 10'h0;
  assign T6406 = T3009[3'h6];
  assign T3013 = T2905 & T6407;
  assign T6407 = {T6408, T3014};
  assign T3014 = ~ T3010;
  assign T6408 = T6409 ? 10'h3ff : 10'h0;
  assign T6409 = T3014[3'h6];
  assign T3015 = T2925 & T3016;
  assign T3016 = 4'ha == T2924;
  assign T3017 = T3022 | T6410;
  assign T6410 = {T6412, T3018};
  assign T3018 = T6411 & T3019;
  assign T3019 = 6'h10;
  assign T6411 = T3020 ? 6'h3f : 6'h0;
  assign T3020 = T3021;
  assign T3021 = 1'h1;
  assign T6412 = T6413 ? 11'h7ff : 11'h0;
  assign T6413 = T3018[3'h5];
  assign T3022 = T2904 & T6414;
  assign T6414 = {T6415, T3023};
  assign T3023 = ~ T3019;
  assign T6415 = T6416 ? 11'h7ff : 11'h0;
  assign T6416 = T3023[3'h5];
  assign T3024 = T2925 & T3025;
  assign T3025 = 4'hb == T2924;
  assign T3026 = T3031 | T6417;
  assign T6417 = {T6419, T3027};
  assign T3027 = T6418 & T3028;
  assign T3028 = 5'h8;
  assign T6418 = T3029 ? 5'h1f : 5'h0;
  assign T3029 = T3030;
  assign T3030 = 1'h1;
  assign T6419 = T6420 ? 12'hfff : 12'h0;
  assign T6420 = T3027[3'h4];
  assign T3031 = T2903 & T6421;
  assign T6421 = {T6422, T3032};
  assign T3032 = ~ T3028;
  assign T6422 = T6423 ? 12'hfff : 12'h0;
  assign T6423 = T3032[3'h4];
  assign T3033 = T2925 & T3034;
  assign T3034 = 4'hc == T2924;
  assign T3035 = T3040 | T6424;
  assign T6424 = {T6426, T3036};
  assign T3036 = T6425 & T3037;
  assign T3037 = 4'h4;
  assign T6425 = T3038 ? 4'hf : 4'h0;
  assign T3038 = T3039;
  assign T3039 = 1'h1;
  assign T6426 = T6427 ? 13'h1fff : 13'h0;
  assign T6427 = T3036[2'h3];
  assign T3040 = T2902 & T6428;
  assign T6428 = {T6429, T3041};
  assign T3041 = ~ T3037;
  assign T6429 = T6430 ? 13'h1fff : 13'h0;
  assign T6430 = T3041[2'h3];
  assign T3042 = T2925 & T3043;
  assign T3043 = 4'hd == T2924;
  assign T3044 = T3049 | T6431;
  assign T6431 = {T6433, T3045};
  assign T3045 = T6432 & T3046;
  assign T3046 = 3'h2;
  assign T6432 = T3047 ? 3'h7 : 3'h0;
  assign T3047 = T3048;
  assign T3048 = 1'h1;
  assign T6433 = T6434 ? 14'h3fff : 14'h0;
  assign T6434 = T3045[2'h2];
  assign T3049 = T2901 & T6435;
  assign T6435 = {T6436, T3050};
  assign T3050 = ~ T3046;
  assign T6436 = T6437 ? 14'h3fff : 14'h0;
  assign T6437 = T3050[2'h2];
  assign T3051 = T2925 & T3052;
  assign T3052 = 4'he == T2924;
  assign T3053 = T3058 | T6438;
  assign T6438 = {T6440, T3054};
  assign T3054 = T6439 & T3055;
  assign T3055 = 2'h1;
  assign T6439 = T3056 ? 2'h3 : 2'h0;
  assign T3056 = T3057;
  assign T3057 = 1'h1;
  assign T6440 = T6441 ? 15'h7fff : 15'h0;
  assign T6441 = T3054[1'h1];
  assign T3058 = T2900 & T6442;
  assign T6442 = {T6443, T3059};
  assign T3059 = ~ T3055;
  assign T6443 = T6444 ? 15'h7fff : 15'h0;
  assign T6444 = T3059[1'h1];
  assign T3060 = T2925 & T3061;
  assign T3061 = 4'hf == T2924;
  assign io_V_wire_en_11 = V_wire_en_11;
  assign V_wire_en_11 = T6445;
  assign T6445 = T3062[4'hf:1'h0];
  assign T3062 = T3223 ? T3216 : T3063;
  assign T3063 = T3214 ? T3207 : T3064;
  assign T3064 = T3205 ? T3198 : T3065;
  assign T3065 = T3196 ? T3189 : T3066;
  assign T3066 = T3187 ? T3180 : T3067;
  assign T3067 = T3178 ? T3171 : T3068;
  assign T3068 = T3169 ? T3162 : T3069;
  assign T3069 = T3160 ? T3153 : T3070;
  assign T3070 = T3151 ? T3144 : T3071;
  assign T3071 = T3142 ? T3135 : T3072;
  assign T3072 = T3133 ? T3126 : T3073;
  assign T3073 = T3124 ? T3117 : T3074;
  assign T3074 = T3115 ? T3108 : T3075;
  assign T3075 = T3106 ? T3099 : T3076;
  assign T3076 = T3097 ? T3090 : T3077;
  assign T3077 = T3085 ? T3078 : 17'h0;
  assign T3078 = T3083 | T3079;
  assign T3079 = T6446 & T3080;
  assign T3080 = 17'h8000;
  assign T6446 = T3081 ? 17'h1ffff : 17'h0;
  assign T3081 = T3082;
  assign T3082 = 1'h1;
  assign T3083 = 17'h0 & T3084;
  assign T3084 = ~ T3080;
  assign T3085 = T3088 & T3086;
  assign T3086 = 4'h0 == T3087;
  assign T3087 = LogicBlockModule_11_io_config_V_out[2'h3:1'h0];
  assign T3088 = T3089;
  assign T3089 = LogicBlockModule_11_io_config_V_out[3'h4];
  assign T3090 = T3095 | T6447;
  assign T6447 = {T6449, T3091};
  assign T3091 = T6448 & T3092;
  assign T3092 = 16'h4000;
  assign T6448 = T3093 ? 16'hffff : 16'h0;
  assign T3093 = T3094;
  assign T3094 = 1'h1;
  assign T6449 = T3091[4'hf];
  assign T3095 = T3077 & T6450;
  assign T6450 = {T6451, T3096};
  assign T3096 = ~ T3092;
  assign T6451 = T3096[4'hf];
  assign T3097 = T3088 & T3098;
  assign T3098 = 4'h1 == T3087;
  assign T3099 = T3104 | T6452;
  assign T6452 = {T6454, T3100};
  assign T3100 = T6453 & T3101;
  assign T3101 = 15'h2000;
  assign T6453 = T3102 ? 15'h7fff : 15'h0;
  assign T3102 = T3103;
  assign T3103 = 1'h1;
  assign T6454 = T6455 ? 2'h3 : 2'h0;
  assign T6455 = T3100[4'he];
  assign T3104 = T3076 & T6456;
  assign T6456 = {T6457, T3105};
  assign T3105 = ~ T3101;
  assign T6457 = T6458 ? 2'h3 : 2'h0;
  assign T6458 = T3105[4'he];
  assign T3106 = T3088 & T3107;
  assign T3107 = 4'h2 == T3087;
  assign T3108 = T3113 | T6459;
  assign T6459 = {T6461, T3109};
  assign T3109 = T6460 & T3110;
  assign T3110 = 14'h1000;
  assign T6460 = T3111 ? 14'h3fff : 14'h0;
  assign T3111 = T3112;
  assign T3112 = 1'h1;
  assign T6461 = T6462 ? 3'h7 : 3'h0;
  assign T6462 = T3109[4'hd];
  assign T3113 = T3075 & T6463;
  assign T6463 = {T6464, T3114};
  assign T3114 = ~ T3110;
  assign T6464 = T6465 ? 3'h7 : 3'h0;
  assign T6465 = T3114[4'hd];
  assign T3115 = T3088 & T3116;
  assign T3116 = 4'h3 == T3087;
  assign T3117 = T3122 | T6466;
  assign T6466 = {T6468, T3118};
  assign T3118 = T6467 & T3119;
  assign T3119 = 13'h800;
  assign T6467 = T3120 ? 13'h1fff : 13'h0;
  assign T3120 = T3121;
  assign T3121 = 1'h1;
  assign T6468 = T6469 ? 4'hf : 4'h0;
  assign T6469 = T3118[4'hc];
  assign T3122 = T3074 & T6470;
  assign T6470 = {T6471, T3123};
  assign T3123 = ~ T3119;
  assign T6471 = T6472 ? 4'hf : 4'h0;
  assign T6472 = T3123[4'hc];
  assign T3124 = T3088 & T3125;
  assign T3125 = 4'h4 == T3087;
  assign T3126 = T3131 | T6473;
  assign T6473 = {T6475, T3127};
  assign T3127 = T6474 & T3128;
  assign T3128 = 12'h400;
  assign T6474 = T3129 ? 12'hfff : 12'h0;
  assign T3129 = T3130;
  assign T3130 = 1'h1;
  assign T6475 = T6476 ? 5'h1f : 5'h0;
  assign T6476 = T3127[4'hb];
  assign T3131 = T3073 & T6477;
  assign T6477 = {T6478, T3132};
  assign T3132 = ~ T3128;
  assign T6478 = T6479 ? 5'h1f : 5'h0;
  assign T6479 = T3132[4'hb];
  assign T3133 = T3088 & T3134;
  assign T3134 = 4'h5 == T3087;
  assign T3135 = T3140 | T6480;
  assign T6480 = {T6482, T3136};
  assign T3136 = T6481 & T3137;
  assign T3137 = 11'h200;
  assign T6481 = T3138 ? 11'h7ff : 11'h0;
  assign T3138 = T3139;
  assign T3139 = 1'h1;
  assign T6482 = T6483 ? 6'h3f : 6'h0;
  assign T6483 = T3136[4'ha];
  assign T3140 = T3072 & T6484;
  assign T6484 = {T6485, T3141};
  assign T3141 = ~ T3137;
  assign T6485 = T6486 ? 6'h3f : 6'h0;
  assign T6486 = T3141[4'ha];
  assign T3142 = T3088 & T3143;
  assign T3143 = 4'h6 == T3087;
  assign T3144 = T3149 | T6487;
  assign T6487 = {T6489, T3145};
  assign T3145 = T6488 & T3146;
  assign T3146 = 10'h100;
  assign T6488 = T3147 ? 10'h3ff : 10'h0;
  assign T3147 = T3148;
  assign T3148 = 1'h1;
  assign T6489 = T6490 ? 7'h7f : 7'h0;
  assign T6490 = T3145[4'h9];
  assign T3149 = T3071 & T6491;
  assign T6491 = {T6492, T3150};
  assign T3150 = ~ T3146;
  assign T6492 = T6493 ? 7'h7f : 7'h0;
  assign T6493 = T3150[4'h9];
  assign T3151 = T3088 & T3152;
  assign T3152 = 4'h7 == T3087;
  assign T3153 = T3158 | T6494;
  assign T6494 = {T6496, T3154};
  assign T3154 = T6495 & T3155;
  assign T3155 = 9'h80;
  assign T6495 = T3156 ? 9'h1ff : 9'h0;
  assign T3156 = T3157;
  assign T3157 = 1'h1;
  assign T6496 = T6497 ? 8'hff : 8'h0;
  assign T6497 = T3154[4'h8];
  assign T3158 = T3070 & T6498;
  assign T6498 = {T6499, T3159};
  assign T3159 = ~ T3155;
  assign T6499 = T6500 ? 8'hff : 8'h0;
  assign T6500 = T3159[4'h8];
  assign T3160 = T3088 & T3161;
  assign T3161 = 4'h8 == T3087;
  assign T3162 = T3167 | T6501;
  assign T6501 = {T6503, T3163};
  assign T3163 = T6502 & T3164;
  assign T3164 = 8'h40;
  assign T6502 = T3165 ? 8'hff : 8'h0;
  assign T3165 = T3166;
  assign T3166 = 1'h1;
  assign T6503 = T6504 ? 9'h1ff : 9'h0;
  assign T6504 = T3163[3'h7];
  assign T3167 = T3069 & T6505;
  assign T6505 = {T6506, T3168};
  assign T3168 = ~ T3164;
  assign T6506 = T6507 ? 9'h1ff : 9'h0;
  assign T6507 = T3168[3'h7];
  assign T3169 = T3088 & T3170;
  assign T3170 = 4'h9 == T3087;
  assign T3171 = T3176 | T6508;
  assign T6508 = {T6510, T3172};
  assign T3172 = T6509 & T3173;
  assign T3173 = 7'h20;
  assign T6509 = T3174 ? 7'h7f : 7'h0;
  assign T3174 = T3175;
  assign T3175 = 1'h1;
  assign T6510 = T6511 ? 10'h3ff : 10'h0;
  assign T6511 = T3172[3'h6];
  assign T3176 = T3068 & T6512;
  assign T6512 = {T6513, T3177};
  assign T3177 = ~ T3173;
  assign T6513 = T6514 ? 10'h3ff : 10'h0;
  assign T6514 = T3177[3'h6];
  assign T3178 = T3088 & T3179;
  assign T3179 = 4'ha == T3087;
  assign T3180 = T3185 | T6515;
  assign T6515 = {T6517, T3181};
  assign T3181 = T6516 & T3182;
  assign T3182 = 6'h10;
  assign T6516 = T3183 ? 6'h3f : 6'h0;
  assign T3183 = T3184;
  assign T3184 = 1'h1;
  assign T6517 = T6518 ? 11'h7ff : 11'h0;
  assign T6518 = T3181[3'h5];
  assign T3185 = T3067 & T6519;
  assign T6519 = {T6520, T3186};
  assign T3186 = ~ T3182;
  assign T6520 = T6521 ? 11'h7ff : 11'h0;
  assign T6521 = T3186[3'h5];
  assign T3187 = T3088 & T3188;
  assign T3188 = 4'hb == T3087;
  assign T3189 = T3194 | T6522;
  assign T6522 = {T6524, T3190};
  assign T3190 = T6523 & T3191;
  assign T3191 = 5'h8;
  assign T6523 = T3192 ? 5'h1f : 5'h0;
  assign T3192 = T3193;
  assign T3193 = 1'h1;
  assign T6524 = T6525 ? 12'hfff : 12'h0;
  assign T6525 = T3190[3'h4];
  assign T3194 = T3066 & T6526;
  assign T6526 = {T6527, T3195};
  assign T3195 = ~ T3191;
  assign T6527 = T6528 ? 12'hfff : 12'h0;
  assign T6528 = T3195[3'h4];
  assign T3196 = T3088 & T3197;
  assign T3197 = 4'hc == T3087;
  assign T3198 = T3203 | T6529;
  assign T6529 = {T6531, T3199};
  assign T3199 = T6530 & T3200;
  assign T3200 = 4'h4;
  assign T6530 = T3201 ? 4'hf : 4'h0;
  assign T3201 = T3202;
  assign T3202 = 1'h1;
  assign T6531 = T6532 ? 13'h1fff : 13'h0;
  assign T6532 = T3199[2'h3];
  assign T3203 = T3065 & T6533;
  assign T6533 = {T6534, T3204};
  assign T3204 = ~ T3200;
  assign T6534 = T6535 ? 13'h1fff : 13'h0;
  assign T6535 = T3204[2'h3];
  assign T3205 = T3088 & T3206;
  assign T3206 = 4'hd == T3087;
  assign T3207 = T3212 | T6536;
  assign T6536 = {T6538, T3208};
  assign T3208 = T6537 & T3209;
  assign T3209 = 3'h2;
  assign T6537 = T3210 ? 3'h7 : 3'h0;
  assign T3210 = T3211;
  assign T3211 = 1'h1;
  assign T6538 = T6539 ? 14'h3fff : 14'h0;
  assign T6539 = T3208[2'h2];
  assign T3212 = T3064 & T6540;
  assign T6540 = {T6541, T3213};
  assign T3213 = ~ T3209;
  assign T6541 = T6542 ? 14'h3fff : 14'h0;
  assign T6542 = T3213[2'h2];
  assign T3214 = T3088 & T3215;
  assign T3215 = 4'he == T3087;
  assign T3216 = T3221 | T6543;
  assign T6543 = {T6545, T3217};
  assign T3217 = T6544 & T3218;
  assign T3218 = 2'h1;
  assign T6544 = T3219 ? 2'h3 : 2'h0;
  assign T3219 = T3220;
  assign T3220 = 1'h1;
  assign T6545 = T6546 ? 15'h7fff : 15'h0;
  assign T6546 = T3217[1'h1];
  assign T3221 = T3063 & T6547;
  assign T6547 = {T6548, T3222};
  assign T3222 = ~ T3218;
  assign T6548 = T6549 ? 15'h7fff : 15'h0;
  assign T6549 = T3222[1'h1];
  assign T3223 = T3088 & T3224;
  assign T3224 = 4'hf == T3087;
  assign io_V_wire_en_12 = V_wire_en_12;
  assign V_wire_en_12 = T6550;
  assign T6550 = T3225[4'hf:1'h0];
  assign T3225 = T3386 ? T3379 : T3226;
  assign T3226 = T3377 ? T3370 : T3227;
  assign T3227 = T3368 ? T3361 : T3228;
  assign T3228 = T3359 ? T3352 : T3229;
  assign T3229 = T3350 ? T3343 : T3230;
  assign T3230 = T3341 ? T3334 : T3231;
  assign T3231 = T3332 ? T3325 : T3232;
  assign T3232 = T3323 ? T3316 : T3233;
  assign T3233 = T3314 ? T3307 : T3234;
  assign T3234 = T3305 ? T3298 : T3235;
  assign T3235 = T3296 ? T3289 : T3236;
  assign T3236 = T3287 ? T3280 : T3237;
  assign T3237 = T3278 ? T3271 : T3238;
  assign T3238 = T3269 ? T3262 : T3239;
  assign T3239 = T3260 ? T3253 : T3240;
  assign T3240 = T3248 ? T3241 : 17'h0;
  assign T3241 = T3246 | T3242;
  assign T3242 = T6551 & T3243;
  assign T3243 = 17'h8000;
  assign T6551 = T3244 ? 17'h1ffff : 17'h0;
  assign T3244 = T3245;
  assign T3245 = 1'h1;
  assign T3246 = 17'h0 & T3247;
  assign T3247 = ~ T3243;
  assign T3248 = T3251 & T3249;
  assign T3249 = 4'h0 == T3250;
  assign T3250 = LogicBlockModule_12_io_config_V_out[2'h3:1'h0];
  assign T3251 = T3252;
  assign T3252 = LogicBlockModule_12_io_config_V_out[3'h4];
  assign T3253 = T3258 | T6552;
  assign T6552 = {T6554, T3254};
  assign T3254 = T6553 & T3255;
  assign T3255 = 16'h4000;
  assign T6553 = T3256 ? 16'hffff : 16'h0;
  assign T3256 = T3257;
  assign T3257 = 1'h1;
  assign T6554 = T3254[4'hf];
  assign T3258 = T3240 & T6555;
  assign T6555 = {T6556, T3259};
  assign T3259 = ~ T3255;
  assign T6556 = T3259[4'hf];
  assign T3260 = T3251 & T3261;
  assign T3261 = 4'h1 == T3250;
  assign T3262 = T3267 | T6557;
  assign T6557 = {T6559, T3263};
  assign T3263 = T6558 & T3264;
  assign T3264 = 15'h2000;
  assign T6558 = T3265 ? 15'h7fff : 15'h0;
  assign T3265 = T3266;
  assign T3266 = 1'h1;
  assign T6559 = T6560 ? 2'h3 : 2'h0;
  assign T6560 = T3263[4'he];
  assign T3267 = T3239 & T6561;
  assign T6561 = {T6562, T3268};
  assign T3268 = ~ T3264;
  assign T6562 = T6563 ? 2'h3 : 2'h0;
  assign T6563 = T3268[4'he];
  assign T3269 = T3251 & T3270;
  assign T3270 = 4'h2 == T3250;
  assign T3271 = T3276 | T6564;
  assign T6564 = {T6566, T3272};
  assign T3272 = T6565 & T3273;
  assign T3273 = 14'h1000;
  assign T6565 = T3274 ? 14'h3fff : 14'h0;
  assign T3274 = T3275;
  assign T3275 = 1'h1;
  assign T6566 = T6567 ? 3'h7 : 3'h0;
  assign T6567 = T3272[4'hd];
  assign T3276 = T3238 & T6568;
  assign T6568 = {T6569, T3277};
  assign T3277 = ~ T3273;
  assign T6569 = T6570 ? 3'h7 : 3'h0;
  assign T6570 = T3277[4'hd];
  assign T3278 = T3251 & T3279;
  assign T3279 = 4'h3 == T3250;
  assign T3280 = T3285 | T6571;
  assign T6571 = {T6573, T3281};
  assign T3281 = T6572 & T3282;
  assign T3282 = 13'h800;
  assign T6572 = T3283 ? 13'h1fff : 13'h0;
  assign T3283 = T3284;
  assign T3284 = 1'h1;
  assign T6573 = T6574 ? 4'hf : 4'h0;
  assign T6574 = T3281[4'hc];
  assign T3285 = T3237 & T6575;
  assign T6575 = {T6576, T3286};
  assign T3286 = ~ T3282;
  assign T6576 = T6577 ? 4'hf : 4'h0;
  assign T6577 = T3286[4'hc];
  assign T3287 = T3251 & T3288;
  assign T3288 = 4'h4 == T3250;
  assign T3289 = T3294 | T6578;
  assign T6578 = {T6580, T3290};
  assign T3290 = T6579 & T3291;
  assign T3291 = 12'h400;
  assign T6579 = T3292 ? 12'hfff : 12'h0;
  assign T3292 = T3293;
  assign T3293 = 1'h1;
  assign T6580 = T6581 ? 5'h1f : 5'h0;
  assign T6581 = T3290[4'hb];
  assign T3294 = T3236 & T6582;
  assign T6582 = {T6583, T3295};
  assign T3295 = ~ T3291;
  assign T6583 = T6584 ? 5'h1f : 5'h0;
  assign T6584 = T3295[4'hb];
  assign T3296 = T3251 & T3297;
  assign T3297 = 4'h5 == T3250;
  assign T3298 = T3303 | T6585;
  assign T6585 = {T6587, T3299};
  assign T3299 = T6586 & T3300;
  assign T3300 = 11'h200;
  assign T6586 = T3301 ? 11'h7ff : 11'h0;
  assign T3301 = T3302;
  assign T3302 = 1'h1;
  assign T6587 = T6588 ? 6'h3f : 6'h0;
  assign T6588 = T3299[4'ha];
  assign T3303 = T3235 & T6589;
  assign T6589 = {T6590, T3304};
  assign T3304 = ~ T3300;
  assign T6590 = T6591 ? 6'h3f : 6'h0;
  assign T6591 = T3304[4'ha];
  assign T3305 = T3251 & T3306;
  assign T3306 = 4'h6 == T3250;
  assign T3307 = T3312 | T6592;
  assign T6592 = {T6594, T3308};
  assign T3308 = T6593 & T3309;
  assign T3309 = 10'h100;
  assign T6593 = T3310 ? 10'h3ff : 10'h0;
  assign T3310 = T3311;
  assign T3311 = 1'h1;
  assign T6594 = T6595 ? 7'h7f : 7'h0;
  assign T6595 = T3308[4'h9];
  assign T3312 = T3234 & T6596;
  assign T6596 = {T6597, T3313};
  assign T3313 = ~ T3309;
  assign T6597 = T6598 ? 7'h7f : 7'h0;
  assign T6598 = T3313[4'h9];
  assign T3314 = T3251 & T3315;
  assign T3315 = 4'h7 == T3250;
  assign T3316 = T3321 | T6599;
  assign T6599 = {T6601, T3317};
  assign T3317 = T6600 & T3318;
  assign T3318 = 9'h80;
  assign T6600 = T3319 ? 9'h1ff : 9'h0;
  assign T3319 = T3320;
  assign T3320 = 1'h1;
  assign T6601 = T6602 ? 8'hff : 8'h0;
  assign T6602 = T3317[4'h8];
  assign T3321 = T3233 & T6603;
  assign T6603 = {T6604, T3322};
  assign T3322 = ~ T3318;
  assign T6604 = T6605 ? 8'hff : 8'h0;
  assign T6605 = T3322[4'h8];
  assign T3323 = T3251 & T3324;
  assign T3324 = 4'h8 == T3250;
  assign T3325 = T3330 | T6606;
  assign T6606 = {T6608, T3326};
  assign T3326 = T6607 & T3327;
  assign T3327 = 8'h40;
  assign T6607 = T3328 ? 8'hff : 8'h0;
  assign T3328 = T3329;
  assign T3329 = 1'h1;
  assign T6608 = T6609 ? 9'h1ff : 9'h0;
  assign T6609 = T3326[3'h7];
  assign T3330 = T3232 & T6610;
  assign T6610 = {T6611, T3331};
  assign T3331 = ~ T3327;
  assign T6611 = T6612 ? 9'h1ff : 9'h0;
  assign T6612 = T3331[3'h7];
  assign T3332 = T3251 & T3333;
  assign T3333 = 4'h9 == T3250;
  assign T3334 = T3339 | T6613;
  assign T6613 = {T6615, T3335};
  assign T3335 = T6614 & T3336;
  assign T3336 = 7'h20;
  assign T6614 = T3337 ? 7'h7f : 7'h0;
  assign T3337 = T3338;
  assign T3338 = 1'h1;
  assign T6615 = T6616 ? 10'h3ff : 10'h0;
  assign T6616 = T3335[3'h6];
  assign T3339 = T3231 & T6617;
  assign T6617 = {T6618, T3340};
  assign T3340 = ~ T3336;
  assign T6618 = T6619 ? 10'h3ff : 10'h0;
  assign T6619 = T3340[3'h6];
  assign T3341 = T3251 & T3342;
  assign T3342 = 4'ha == T3250;
  assign T3343 = T3348 | T6620;
  assign T6620 = {T6622, T3344};
  assign T3344 = T6621 & T3345;
  assign T3345 = 6'h10;
  assign T6621 = T3346 ? 6'h3f : 6'h0;
  assign T3346 = T3347;
  assign T3347 = 1'h1;
  assign T6622 = T6623 ? 11'h7ff : 11'h0;
  assign T6623 = T3344[3'h5];
  assign T3348 = T3230 & T6624;
  assign T6624 = {T6625, T3349};
  assign T3349 = ~ T3345;
  assign T6625 = T6626 ? 11'h7ff : 11'h0;
  assign T6626 = T3349[3'h5];
  assign T3350 = T3251 & T3351;
  assign T3351 = 4'hb == T3250;
  assign T3352 = T3357 | T6627;
  assign T6627 = {T6629, T3353};
  assign T3353 = T6628 & T3354;
  assign T3354 = 5'h8;
  assign T6628 = T3355 ? 5'h1f : 5'h0;
  assign T3355 = T3356;
  assign T3356 = 1'h1;
  assign T6629 = T6630 ? 12'hfff : 12'h0;
  assign T6630 = T3353[3'h4];
  assign T3357 = T3229 & T6631;
  assign T6631 = {T6632, T3358};
  assign T3358 = ~ T3354;
  assign T6632 = T6633 ? 12'hfff : 12'h0;
  assign T6633 = T3358[3'h4];
  assign T3359 = T3251 & T3360;
  assign T3360 = 4'hc == T3250;
  assign T3361 = T3366 | T6634;
  assign T6634 = {T6636, T3362};
  assign T3362 = T6635 & T3363;
  assign T3363 = 4'h4;
  assign T6635 = T3364 ? 4'hf : 4'h0;
  assign T3364 = T3365;
  assign T3365 = 1'h1;
  assign T6636 = T6637 ? 13'h1fff : 13'h0;
  assign T6637 = T3362[2'h3];
  assign T3366 = T3228 & T6638;
  assign T6638 = {T6639, T3367};
  assign T3367 = ~ T3363;
  assign T6639 = T6640 ? 13'h1fff : 13'h0;
  assign T6640 = T3367[2'h3];
  assign T3368 = T3251 & T3369;
  assign T3369 = 4'hd == T3250;
  assign T3370 = T3375 | T6641;
  assign T6641 = {T6643, T3371};
  assign T3371 = T6642 & T3372;
  assign T3372 = 3'h2;
  assign T6642 = T3373 ? 3'h7 : 3'h0;
  assign T3373 = T3374;
  assign T3374 = 1'h1;
  assign T6643 = T6644 ? 14'h3fff : 14'h0;
  assign T6644 = T3371[2'h2];
  assign T3375 = T3227 & T6645;
  assign T6645 = {T6646, T3376};
  assign T3376 = ~ T3372;
  assign T6646 = T6647 ? 14'h3fff : 14'h0;
  assign T6647 = T3376[2'h2];
  assign T3377 = T3251 & T3378;
  assign T3378 = 4'he == T3250;
  assign T3379 = T3384 | T6648;
  assign T6648 = {T6650, T3380};
  assign T3380 = T6649 & T3381;
  assign T3381 = 2'h1;
  assign T6649 = T3382 ? 2'h3 : 2'h0;
  assign T3382 = T3383;
  assign T3383 = 1'h1;
  assign T6650 = T6651 ? 15'h7fff : 15'h0;
  assign T6651 = T3380[1'h1];
  assign T3384 = T3226 & T6652;
  assign T6652 = {T6653, T3385};
  assign T3385 = ~ T3381;
  assign T6653 = T6654 ? 15'h7fff : 15'h0;
  assign T6654 = T3385[1'h1];
  assign T3386 = T3251 & T3387;
  assign T3387 = 4'hf == T3250;
  assign io_V_wire_en_13 = V_wire_en_13;
  assign V_wire_en_13 = T6655;
  assign T6655 = T3388[4'hf:1'h0];
  assign T3388 = T3549 ? T3542 : T3389;
  assign T3389 = T3540 ? T3533 : T3390;
  assign T3390 = T3531 ? T3524 : T3391;
  assign T3391 = T3522 ? T3515 : T3392;
  assign T3392 = T3513 ? T3506 : T3393;
  assign T3393 = T3504 ? T3497 : T3394;
  assign T3394 = T3495 ? T3488 : T3395;
  assign T3395 = T3486 ? T3479 : T3396;
  assign T3396 = T3477 ? T3470 : T3397;
  assign T3397 = T3468 ? T3461 : T3398;
  assign T3398 = T3459 ? T3452 : T3399;
  assign T3399 = T3450 ? T3443 : T3400;
  assign T3400 = T3441 ? T3434 : T3401;
  assign T3401 = T3432 ? T3425 : T3402;
  assign T3402 = T3423 ? T3416 : T3403;
  assign T3403 = T3411 ? T3404 : 17'h0;
  assign T3404 = T3409 | T3405;
  assign T3405 = T6656 & T3406;
  assign T3406 = 17'h8000;
  assign T6656 = T3407 ? 17'h1ffff : 17'h0;
  assign T3407 = T3408;
  assign T3408 = 1'h1;
  assign T3409 = 17'h0 & T3410;
  assign T3410 = ~ T3406;
  assign T3411 = T3414 & T3412;
  assign T3412 = 4'h0 == T3413;
  assign T3413 = LogicBlockModule_13_io_config_V_out[2'h3:1'h0];
  assign T3414 = T3415;
  assign T3415 = LogicBlockModule_13_io_config_V_out[3'h4];
  assign T3416 = T3421 | T6657;
  assign T6657 = {T6659, T3417};
  assign T3417 = T6658 & T3418;
  assign T3418 = 16'h4000;
  assign T6658 = T3419 ? 16'hffff : 16'h0;
  assign T3419 = T3420;
  assign T3420 = 1'h1;
  assign T6659 = T3417[4'hf];
  assign T3421 = T3403 & T6660;
  assign T6660 = {T6661, T3422};
  assign T3422 = ~ T3418;
  assign T6661 = T3422[4'hf];
  assign T3423 = T3414 & T3424;
  assign T3424 = 4'h1 == T3413;
  assign T3425 = T3430 | T6662;
  assign T6662 = {T6664, T3426};
  assign T3426 = T6663 & T3427;
  assign T3427 = 15'h2000;
  assign T6663 = T3428 ? 15'h7fff : 15'h0;
  assign T3428 = T3429;
  assign T3429 = 1'h1;
  assign T6664 = T6665 ? 2'h3 : 2'h0;
  assign T6665 = T3426[4'he];
  assign T3430 = T3402 & T6666;
  assign T6666 = {T6667, T3431};
  assign T3431 = ~ T3427;
  assign T6667 = T6668 ? 2'h3 : 2'h0;
  assign T6668 = T3431[4'he];
  assign T3432 = T3414 & T3433;
  assign T3433 = 4'h2 == T3413;
  assign T3434 = T3439 | T6669;
  assign T6669 = {T6671, T3435};
  assign T3435 = T6670 & T3436;
  assign T3436 = 14'h1000;
  assign T6670 = T3437 ? 14'h3fff : 14'h0;
  assign T3437 = T3438;
  assign T3438 = 1'h1;
  assign T6671 = T6672 ? 3'h7 : 3'h0;
  assign T6672 = T3435[4'hd];
  assign T3439 = T3401 & T6673;
  assign T6673 = {T6674, T3440};
  assign T3440 = ~ T3436;
  assign T6674 = T6675 ? 3'h7 : 3'h0;
  assign T6675 = T3440[4'hd];
  assign T3441 = T3414 & T3442;
  assign T3442 = 4'h3 == T3413;
  assign T3443 = T3448 | T6676;
  assign T6676 = {T6678, T3444};
  assign T3444 = T6677 & T3445;
  assign T3445 = 13'h800;
  assign T6677 = T3446 ? 13'h1fff : 13'h0;
  assign T3446 = T3447;
  assign T3447 = 1'h1;
  assign T6678 = T6679 ? 4'hf : 4'h0;
  assign T6679 = T3444[4'hc];
  assign T3448 = T3400 & T6680;
  assign T6680 = {T6681, T3449};
  assign T3449 = ~ T3445;
  assign T6681 = T6682 ? 4'hf : 4'h0;
  assign T6682 = T3449[4'hc];
  assign T3450 = T3414 & T3451;
  assign T3451 = 4'h4 == T3413;
  assign T3452 = T3457 | T6683;
  assign T6683 = {T6685, T3453};
  assign T3453 = T6684 & T3454;
  assign T3454 = 12'h400;
  assign T6684 = T3455 ? 12'hfff : 12'h0;
  assign T3455 = T3456;
  assign T3456 = 1'h1;
  assign T6685 = T6686 ? 5'h1f : 5'h0;
  assign T6686 = T3453[4'hb];
  assign T3457 = T3399 & T6687;
  assign T6687 = {T6688, T3458};
  assign T3458 = ~ T3454;
  assign T6688 = T6689 ? 5'h1f : 5'h0;
  assign T6689 = T3458[4'hb];
  assign T3459 = T3414 & T3460;
  assign T3460 = 4'h5 == T3413;
  assign T3461 = T3466 | T6690;
  assign T6690 = {T6692, T3462};
  assign T3462 = T6691 & T3463;
  assign T3463 = 11'h200;
  assign T6691 = T3464 ? 11'h7ff : 11'h0;
  assign T3464 = T3465;
  assign T3465 = 1'h1;
  assign T6692 = T6693 ? 6'h3f : 6'h0;
  assign T6693 = T3462[4'ha];
  assign T3466 = T3398 & T6694;
  assign T6694 = {T6695, T3467};
  assign T3467 = ~ T3463;
  assign T6695 = T6696 ? 6'h3f : 6'h0;
  assign T6696 = T3467[4'ha];
  assign T3468 = T3414 & T3469;
  assign T3469 = 4'h6 == T3413;
  assign T3470 = T3475 | T6697;
  assign T6697 = {T6699, T3471};
  assign T3471 = T6698 & T3472;
  assign T3472 = 10'h100;
  assign T6698 = T3473 ? 10'h3ff : 10'h0;
  assign T3473 = T3474;
  assign T3474 = 1'h1;
  assign T6699 = T6700 ? 7'h7f : 7'h0;
  assign T6700 = T3471[4'h9];
  assign T3475 = T3397 & T6701;
  assign T6701 = {T6702, T3476};
  assign T3476 = ~ T3472;
  assign T6702 = T6703 ? 7'h7f : 7'h0;
  assign T6703 = T3476[4'h9];
  assign T3477 = T3414 & T3478;
  assign T3478 = 4'h7 == T3413;
  assign T3479 = T3484 | T6704;
  assign T6704 = {T6706, T3480};
  assign T3480 = T6705 & T3481;
  assign T3481 = 9'h80;
  assign T6705 = T3482 ? 9'h1ff : 9'h0;
  assign T3482 = T3483;
  assign T3483 = 1'h1;
  assign T6706 = T6707 ? 8'hff : 8'h0;
  assign T6707 = T3480[4'h8];
  assign T3484 = T3396 & T6708;
  assign T6708 = {T6709, T3485};
  assign T3485 = ~ T3481;
  assign T6709 = T6710 ? 8'hff : 8'h0;
  assign T6710 = T3485[4'h8];
  assign T3486 = T3414 & T3487;
  assign T3487 = 4'h8 == T3413;
  assign T3488 = T3493 | T6711;
  assign T6711 = {T6713, T3489};
  assign T3489 = T6712 & T3490;
  assign T3490 = 8'h40;
  assign T6712 = T3491 ? 8'hff : 8'h0;
  assign T3491 = T3492;
  assign T3492 = 1'h1;
  assign T6713 = T6714 ? 9'h1ff : 9'h0;
  assign T6714 = T3489[3'h7];
  assign T3493 = T3395 & T6715;
  assign T6715 = {T6716, T3494};
  assign T3494 = ~ T3490;
  assign T6716 = T6717 ? 9'h1ff : 9'h0;
  assign T6717 = T3494[3'h7];
  assign T3495 = T3414 & T3496;
  assign T3496 = 4'h9 == T3413;
  assign T3497 = T3502 | T6718;
  assign T6718 = {T6720, T3498};
  assign T3498 = T6719 & T3499;
  assign T3499 = 7'h20;
  assign T6719 = T3500 ? 7'h7f : 7'h0;
  assign T3500 = T3501;
  assign T3501 = 1'h1;
  assign T6720 = T6721 ? 10'h3ff : 10'h0;
  assign T6721 = T3498[3'h6];
  assign T3502 = T3394 & T6722;
  assign T6722 = {T6723, T3503};
  assign T3503 = ~ T3499;
  assign T6723 = T6724 ? 10'h3ff : 10'h0;
  assign T6724 = T3503[3'h6];
  assign T3504 = T3414 & T3505;
  assign T3505 = 4'ha == T3413;
  assign T3506 = T3511 | T6725;
  assign T6725 = {T6727, T3507};
  assign T3507 = T6726 & T3508;
  assign T3508 = 6'h10;
  assign T6726 = T3509 ? 6'h3f : 6'h0;
  assign T3509 = T3510;
  assign T3510 = 1'h1;
  assign T6727 = T6728 ? 11'h7ff : 11'h0;
  assign T6728 = T3507[3'h5];
  assign T3511 = T3393 & T6729;
  assign T6729 = {T6730, T3512};
  assign T3512 = ~ T3508;
  assign T6730 = T6731 ? 11'h7ff : 11'h0;
  assign T6731 = T3512[3'h5];
  assign T3513 = T3414 & T3514;
  assign T3514 = 4'hb == T3413;
  assign T3515 = T3520 | T6732;
  assign T6732 = {T6734, T3516};
  assign T3516 = T6733 & T3517;
  assign T3517 = 5'h8;
  assign T6733 = T3518 ? 5'h1f : 5'h0;
  assign T3518 = T3519;
  assign T3519 = 1'h1;
  assign T6734 = T6735 ? 12'hfff : 12'h0;
  assign T6735 = T3516[3'h4];
  assign T3520 = T3392 & T6736;
  assign T6736 = {T6737, T3521};
  assign T3521 = ~ T3517;
  assign T6737 = T6738 ? 12'hfff : 12'h0;
  assign T6738 = T3521[3'h4];
  assign T3522 = T3414 & T3523;
  assign T3523 = 4'hc == T3413;
  assign T3524 = T3529 | T6739;
  assign T6739 = {T6741, T3525};
  assign T3525 = T6740 & T3526;
  assign T3526 = 4'h4;
  assign T6740 = T3527 ? 4'hf : 4'h0;
  assign T3527 = T3528;
  assign T3528 = 1'h1;
  assign T6741 = T6742 ? 13'h1fff : 13'h0;
  assign T6742 = T3525[2'h3];
  assign T3529 = T3391 & T6743;
  assign T6743 = {T6744, T3530};
  assign T3530 = ~ T3526;
  assign T6744 = T6745 ? 13'h1fff : 13'h0;
  assign T6745 = T3530[2'h3];
  assign T3531 = T3414 & T3532;
  assign T3532 = 4'hd == T3413;
  assign T3533 = T3538 | T6746;
  assign T6746 = {T6748, T3534};
  assign T3534 = T6747 & T3535;
  assign T3535 = 3'h2;
  assign T6747 = T3536 ? 3'h7 : 3'h0;
  assign T3536 = T3537;
  assign T3537 = 1'h1;
  assign T6748 = T6749 ? 14'h3fff : 14'h0;
  assign T6749 = T3534[2'h2];
  assign T3538 = T3390 & T6750;
  assign T6750 = {T6751, T3539};
  assign T3539 = ~ T3535;
  assign T6751 = T6752 ? 14'h3fff : 14'h0;
  assign T6752 = T3539[2'h2];
  assign T3540 = T3414 & T3541;
  assign T3541 = 4'he == T3413;
  assign T3542 = T3547 | T6753;
  assign T6753 = {T6755, T3543};
  assign T3543 = T6754 & T3544;
  assign T3544 = 2'h1;
  assign T6754 = T3545 ? 2'h3 : 2'h0;
  assign T3545 = T3546;
  assign T3546 = 1'h1;
  assign T6755 = T6756 ? 15'h7fff : 15'h0;
  assign T6756 = T3543[1'h1];
  assign T3547 = T3389 & T6757;
  assign T6757 = {T6758, T3548};
  assign T3548 = ~ T3544;
  assign T6758 = T6759 ? 15'h7fff : 15'h0;
  assign T6759 = T3548[1'h1];
  assign T3549 = T3414 & T3550;
  assign T3550 = 4'hf == T3413;
  assign io_V_wire_en_14 = V_wire_en_14;
  assign V_wire_en_14 = T6760;
  assign T6760 = T3551[4'hf:1'h0];
  assign T3551 = T3712 ? T3705 : T3552;
  assign T3552 = T3703 ? T3696 : T3553;
  assign T3553 = T3694 ? T3687 : T3554;
  assign T3554 = T3685 ? T3678 : T3555;
  assign T3555 = T3676 ? T3669 : T3556;
  assign T3556 = T3667 ? T3660 : T3557;
  assign T3557 = T3658 ? T3651 : T3558;
  assign T3558 = T3649 ? T3642 : T3559;
  assign T3559 = T3640 ? T3633 : T3560;
  assign T3560 = T3631 ? T3624 : T3561;
  assign T3561 = T3622 ? T3615 : T3562;
  assign T3562 = T3613 ? T3606 : T3563;
  assign T3563 = T3604 ? T3597 : T3564;
  assign T3564 = T3595 ? T3588 : T3565;
  assign T3565 = T3586 ? T3579 : T3566;
  assign T3566 = T3574 ? T3567 : 17'h0;
  assign T3567 = T3572 | T3568;
  assign T3568 = T6761 & T3569;
  assign T3569 = 17'h8000;
  assign T6761 = T3570 ? 17'h1ffff : 17'h0;
  assign T3570 = T3571;
  assign T3571 = 1'h1;
  assign T3572 = 17'h0 & T3573;
  assign T3573 = ~ T3569;
  assign T3574 = T3577 & T3575;
  assign T3575 = 4'h0 == T3576;
  assign T3576 = LogicBlockModule_14_io_config_V_out[2'h3:1'h0];
  assign T3577 = T3578;
  assign T3578 = LogicBlockModule_14_io_config_V_out[3'h4];
  assign T3579 = T3584 | T6762;
  assign T6762 = {T6764, T3580};
  assign T3580 = T6763 & T3581;
  assign T3581 = 16'h4000;
  assign T6763 = T3582 ? 16'hffff : 16'h0;
  assign T3582 = T3583;
  assign T3583 = 1'h1;
  assign T6764 = T3580[4'hf];
  assign T3584 = T3566 & T6765;
  assign T6765 = {T6766, T3585};
  assign T3585 = ~ T3581;
  assign T6766 = T3585[4'hf];
  assign T3586 = T3577 & T3587;
  assign T3587 = 4'h1 == T3576;
  assign T3588 = T3593 | T6767;
  assign T6767 = {T6769, T3589};
  assign T3589 = T6768 & T3590;
  assign T3590 = 15'h2000;
  assign T6768 = T3591 ? 15'h7fff : 15'h0;
  assign T3591 = T3592;
  assign T3592 = 1'h1;
  assign T6769 = T6770 ? 2'h3 : 2'h0;
  assign T6770 = T3589[4'he];
  assign T3593 = T3565 & T6771;
  assign T6771 = {T6772, T3594};
  assign T3594 = ~ T3590;
  assign T6772 = T6773 ? 2'h3 : 2'h0;
  assign T6773 = T3594[4'he];
  assign T3595 = T3577 & T3596;
  assign T3596 = 4'h2 == T3576;
  assign T3597 = T3602 | T6774;
  assign T6774 = {T6776, T3598};
  assign T3598 = T6775 & T3599;
  assign T3599 = 14'h1000;
  assign T6775 = T3600 ? 14'h3fff : 14'h0;
  assign T3600 = T3601;
  assign T3601 = 1'h1;
  assign T6776 = T6777 ? 3'h7 : 3'h0;
  assign T6777 = T3598[4'hd];
  assign T3602 = T3564 & T6778;
  assign T6778 = {T6779, T3603};
  assign T3603 = ~ T3599;
  assign T6779 = T6780 ? 3'h7 : 3'h0;
  assign T6780 = T3603[4'hd];
  assign T3604 = T3577 & T3605;
  assign T3605 = 4'h3 == T3576;
  assign T3606 = T3611 | T6781;
  assign T6781 = {T6783, T3607};
  assign T3607 = T6782 & T3608;
  assign T3608 = 13'h800;
  assign T6782 = T3609 ? 13'h1fff : 13'h0;
  assign T3609 = T3610;
  assign T3610 = 1'h1;
  assign T6783 = T6784 ? 4'hf : 4'h0;
  assign T6784 = T3607[4'hc];
  assign T3611 = T3563 & T6785;
  assign T6785 = {T6786, T3612};
  assign T3612 = ~ T3608;
  assign T6786 = T6787 ? 4'hf : 4'h0;
  assign T6787 = T3612[4'hc];
  assign T3613 = T3577 & T3614;
  assign T3614 = 4'h4 == T3576;
  assign T3615 = T3620 | T6788;
  assign T6788 = {T6790, T3616};
  assign T3616 = T6789 & T3617;
  assign T3617 = 12'h400;
  assign T6789 = T3618 ? 12'hfff : 12'h0;
  assign T3618 = T3619;
  assign T3619 = 1'h1;
  assign T6790 = T6791 ? 5'h1f : 5'h0;
  assign T6791 = T3616[4'hb];
  assign T3620 = T3562 & T6792;
  assign T6792 = {T6793, T3621};
  assign T3621 = ~ T3617;
  assign T6793 = T6794 ? 5'h1f : 5'h0;
  assign T6794 = T3621[4'hb];
  assign T3622 = T3577 & T3623;
  assign T3623 = 4'h5 == T3576;
  assign T3624 = T3629 | T6795;
  assign T6795 = {T6797, T3625};
  assign T3625 = T6796 & T3626;
  assign T3626 = 11'h200;
  assign T6796 = T3627 ? 11'h7ff : 11'h0;
  assign T3627 = T3628;
  assign T3628 = 1'h1;
  assign T6797 = T6798 ? 6'h3f : 6'h0;
  assign T6798 = T3625[4'ha];
  assign T3629 = T3561 & T6799;
  assign T6799 = {T6800, T3630};
  assign T3630 = ~ T3626;
  assign T6800 = T6801 ? 6'h3f : 6'h0;
  assign T6801 = T3630[4'ha];
  assign T3631 = T3577 & T3632;
  assign T3632 = 4'h6 == T3576;
  assign T3633 = T3638 | T6802;
  assign T6802 = {T6804, T3634};
  assign T3634 = T6803 & T3635;
  assign T3635 = 10'h100;
  assign T6803 = T3636 ? 10'h3ff : 10'h0;
  assign T3636 = T3637;
  assign T3637 = 1'h1;
  assign T6804 = T6805 ? 7'h7f : 7'h0;
  assign T6805 = T3634[4'h9];
  assign T3638 = T3560 & T6806;
  assign T6806 = {T6807, T3639};
  assign T3639 = ~ T3635;
  assign T6807 = T6808 ? 7'h7f : 7'h0;
  assign T6808 = T3639[4'h9];
  assign T3640 = T3577 & T3641;
  assign T3641 = 4'h7 == T3576;
  assign T3642 = T3647 | T6809;
  assign T6809 = {T6811, T3643};
  assign T3643 = T6810 & T3644;
  assign T3644 = 9'h80;
  assign T6810 = T3645 ? 9'h1ff : 9'h0;
  assign T3645 = T3646;
  assign T3646 = 1'h1;
  assign T6811 = T6812 ? 8'hff : 8'h0;
  assign T6812 = T3643[4'h8];
  assign T3647 = T3559 & T6813;
  assign T6813 = {T6814, T3648};
  assign T3648 = ~ T3644;
  assign T6814 = T6815 ? 8'hff : 8'h0;
  assign T6815 = T3648[4'h8];
  assign T3649 = T3577 & T3650;
  assign T3650 = 4'h8 == T3576;
  assign T3651 = T3656 | T6816;
  assign T6816 = {T6818, T3652};
  assign T3652 = T6817 & T3653;
  assign T3653 = 8'h40;
  assign T6817 = T3654 ? 8'hff : 8'h0;
  assign T3654 = T3655;
  assign T3655 = 1'h1;
  assign T6818 = T6819 ? 9'h1ff : 9'h0;
  assign T6819 = T3652[3'h7];
  assign T3656 = T3558 & T6820;
  assign T6820 = {T6821, T3657};
  assign T3657 = ~ T3653;
  assign T6821 = T6822 ? 9'h1ff : 9'h0;
  assign T6822 = T3657[3'h7];
  assign T3658 = T3577 & T3659;
  assign T3659 = 4'h9 == T3576;
  assign T3660 = T3665 | T6823;
  assign T6823 = {T6825, T3661};
  assign T3661 = T6824 & T3662;
  assign T3662 = 7'h20;
  assign T6824 = T3663 ? 7'h7f : 7'h0;
  assign T3663 = T3664;
  assign T3664 = 1'h1;
  assign T6825 = T6826 ? 10'h3ff : 10'h0;
  assign T6826 = T3661[3'h6];
  assign T3665 = T3557 & T6827;
  assign T6827 = {T6828, T3666};
  assign T3666 = ~ T3662;
  assign T6828 = T6829 ? 10'h3ff : 10'h0;
  assign T6829 = T3666[3'h6];
  assign T3667 = T3577 & T3668;
  assign T3668 = 4'ha == T3576;
  assign T3669 = T3674 | T6830;
  assign T6830 = {T6832, T3670};
  assign T3670 = T6831 & T3671;
  assign T3671 = 6'h10;
  assign T6831 = T3672 ? 6'h3f : 6'h0;
  assign T3672 = T3673;
  assign T3673 = 1'h1;
  assign T6832 = T6833 ? 11'h7ff : 11'h0;
  assign T6833 = T3670[3'h5];
  assign T3674 = T3556 & T6834;
  assign T6834 = {T6835, T3675};
  assign T3675 = ~ T3671;
  assign T6835 = T6836 ? 11'h7ff : 11'h0;
  assign T6836 = T3675[3'h5];
  assign T3676 = T3577 & T3677;
  assign T3677 = 4'hb == T3576;
  assign T3678 = T3683 | T6837;
  assign T6837 = {T6839, T3679};
  assign T3679 = T6838 & T3680;
  assign T3680 = 5'h8;
  assign T6838 = T3681 ? 5'h1f : 5'h0;
  assign T3681 = T3682;
  assign T3682 = 1'h1;
  assign T6839 = T6840 ? 12'hfff : 12'h0;
  assign T6840 = T3679[3'h4];
  assign T3683 = T3555 & T6841;
  assign T6841 = {T6842, T3684};
  assign T3684 = ~ T3680;
  assign T6842 = T6843 ? 12'hfff : 12'h0;
  assign T6843 = T3684[3'h4];
  assign T3685 = T3577 & T3686;
  assign T3686 = 4'hc == T3576;
  assign T3687 = T3692 | T6844;
  assign T6844 = {T6846, T3688};
  assign T3688 = T6845 & T3689;
  assign T3689 = 4'h4;
  assign T6845 = T3690 ? 4'hf : 4'h0;
  assign T3690 = T3691;
  assign T3691 = 1'h1;
  assign T6846 = T6847 ? 13'h1fff : 13'h0;
  assign T6847 = T3688[2'h3];
  assign T3692 = T3554 & T6848;
  assign T6848 = {T6849, T3693};
  assign T3693 = ~ T3689;
  assign T6849 = T6850 ? 13'h1fff : 13'h0;
  assign T6850 = T3693[2'h3];
  assign T3694 = T3577 & T3695;
  assign T3695 = 4'hd == T3576;
  assign T3696 = T3701 | T6851;
  assign T6851 = {T6853, T3697};
  assign T3697 = T6852 & T3698;
  assign T3698 = 3'h2;
  assign T6852 = T3699 ? 3'h7 : 3'h0;
  assign T3699 = T3700;
  assign T3700 = 1'h1;
  assign T6853 = T6854 ? 14'h3fff : 14'h0;
  assign T6854 = T3697[2'h2];
  assign T3701 = T3553 & T6855;
  assign T6855 = {T6856, T3702};
  assign T3702 = ~ T3698;
  assign T6856 = T6857 ? 14'h3fff : 14'h0;
  assign T6857 = T3702[2'h2];
  assign T3703 = T3577 & T3704;
  assign T3704 = 4'he == T3576;
  assign T3705 = T3710 | T6858;
  assign T6858 = {T6860, T3706};
  assign T3706 = T6859 & T3707;
  assign T3707 = 2'h1;
  assign T6859 = T3708 ? 2'h3 : 2'h0;
  assign T3708 = T3709;
  assign T3709 = 1'h1;
  assign T6860 = T6861 ? 15'h7fff : 15'h0;
  assign T6861 = T3706[1'h1];
  assign T3710 = T3552 & T6862;
  assign T6862 = {T6863, T3711};
  assign T3711 = ~ T3707;
  assign T6863 = T6864 ? 15'h7fff : 15'h0;
  assign T6864 = T3711[1'h1];
  assign T3712 = T3577 & T3713;
  assign T3713 = 4'hf == T3576;
  assign io_V_wire_en_15 = V_wire_en_15;
  assign V_wire_en_15 = T6865;
  assign T6865 = T3714[4'hf:1'h0];
  assign T3714 = T3875 ? T3868 : T3715;
  assign T3715 = T3866 ? T3859 : T3716;
  assign T3716 = T3857 ? T3850 : T3717;
  assign T3717 = T3848 ? T3841 : T3718;
  assign T3718 = T3839 ? T3832 : T3719;
  assign T3719 = T3830 ? T3823 : T3720;
  assign T3720 = T3821 ? T3814 : T3721;
  assign T3721 = T3812 ? T3805 : T3722;
  assign T3722 = T3803 ? T3796 : T3723;
  assign T3723 = T3794 ? T3787 : T3724;
  assign T3724 = T3785 ? T3778 : T3725;
  assign T3725 = T3776 ? T3769 : T3726;
  assign T3726 = T3767 ? T3760 : T3727;
  assign T3727 = T3758 ? T3751 : T3728;
  assign T3728 = T3749 ? T3742 : T3729;
  assign T3729 = T3737 ? T3730 : 17'h0;
  assign T3730 = T3735 | T3731;
  assign T3731 = T6866 & T3732;
  assign T3732 = 17'h8000;
  assign T6866 = T3733 ? 17'h1ffff : 17'h0;
  assign T3733 = T3734;
  assign T3734 = 1'h1;
  assign T3735 = 17'h0 & T3736;
  assign T3736 = ~ T3732;
  assign T3737 = T3740 & T3738;
  assign T3738 = 4'h0 == T3739;
  assign T3739 = LogicBlockModule_15_io_config_V_out[2'h3:1'h0];
  assign T3740 = T3741;
  assign T3741 = LogicBlockModule_15_io_config_V_out[3'h4];
  assign T3742 = T3747 | T6867;
  assign T6867 = {T6869, T3743};
  assign T3743 = T6868 & T3744;
  assign T3744 = 16'h4000;
  assign T6868 = T3745 ? 16'hffff : 16'h0;
  assign T3745 = T3746;
  assign T3746 = 1'h1;
  assign T6869 = T3743[4'hf];
  assign T3747 = T3729 & T6870;
  assign T6870 = {T6871, T3748};
  assign T3748 = ~ T3744;
  assign T6871 = T3748[4'hf];
  assign T3749 = T3740 & T3750;
  assign T3750 = 4'h1 == T3739;
  assign T3751 = T3756 | T6872;
  assign T6872 = {T6874, T3752};
  assign T3752 = T6873 & T3753;
  assign T3753 = 15'h2000;
  assign T6873 = T3754 ? 15'h7fff : 15'h0;
  assign T3754 = T3755;
  assign T3755 = 1'h1;
  assign T6874 = T6875 ? 2'h3 : 2'h0;
  assign T6875 = T3752[4'he];
  assign T3756 = T3728 & T6876;
  assign T6876 = {T6877, T3757};
  assign T3757 = ~ T3753;
  assign T6877 = T6878 ? 2'h3 : 2'h0;
  assign T6878 = T3757[4'he];
  assign T3758 = T3740 & T3759;
  assign T3759 = 4'h2 == T3739;
  assign T3760 = T3765 | T6879;
  assign T6879 = {T6881, T3761};
  assign T3761 = T6880 & T3762;
  assign T3762 = 14'h1000;
  assign T6880 = T3763 ? 14'h3fff : 14'h0;
  assign T3763 = T3764;
  assign T3764 = 1'h1;
  assign T6881 = T6882 ? 3'h7 : 3'h0;
  assign T6882 = T3761[4'hd];
  assign T3765 = T3727 & T6883;
  assign T6883 = {T6884, T3766};
  assign T3766 = ~ T3762;
  assign T6884 = T6885 ? 3'h7 : 3'h0;
  assign T6885 = T3766[4'hd];
  assign T3767 = T3740 & T3768;
  assign T3768 = 4'h3 == T3739;
  assign T3769 = T3774 | T6886;
  assign T6886 = {T6888, T3770};
  assign T3770 = T6887 & T3771;
  assign T3771 = 13'h800;
  assign T6887 = T3772 ? 13'h1fff : 13'h0;
  assign T3772 = T3773;
  assign T3773 = 1'h1;
  assign T6888 = T6889 ? 4'hf : 4'h0;
  assign T6889 = T3770[4'hc];
  assign T3774 = T3726 & T6890;
  assign T6890 = {T6891, T3775};
  assign T3775 = ~ T3771;
  assign T6891 = T6892 ? 4'hf : 4'h0;
  assign T6892 = T3775[4'hc];
  assign T3776 = T3740 & T3777;
  assign T3777 = 4'h4 == T3739;
  assign T3778 = T3783 | T6893;
  assign T6893 = {T6895, T3779};
  assign T3779 = T6894 & T3780;
  assign T3780 = 12'h400;
  assign T6894 = T3781 ? 12'hfff : 12'h0;
  assign T3781 = T3782;
  assign T3782 = 1'h1;
  assign T6895 = T6896 ? 5'h1f : 5'h0;
  assign T6896 = T3779[4'hb];
  assign T3783 = T3725 & T6897;
  assign T6897 = {T6898, T3784};
  assign T3784 = ~ T3780;
  assign T6898 = T6899 ? 5'h1f : 5'h0;
  assign T6899 = T3784[4'hb];
  assign T3785 = T3740 & T3786;
  assign T3786 = 4'h5 == T3739;
  assign T3787 = T3792 | T6900;
  assign T6900 = {T6902, T3788};
  assign T3788 = T6901 & T3789;
  assign T3789 = 11'h200;
  assign T6901 = T3790 ? 11'h7ff : 11'h0;
  assign T3790 = T3791;
  assign T3791 = 1'h1;
  assign T6902 = T6903 ? 6'h3f : 6'h0;
  assign T6903 = T3788[4'ha];
  assign T3792 = T3724 & T6904;
  assign T6904 = {T6905, T3793};
  assign T3793 = ~ T3789;
  assign T6905 = T6906 ? 6'h3f : 6'h0;
  assign T6906 = T3793[4'ha];
  assign T3794 = T3740 & T3795;
  assign T3795 = 4'h6 == T3739;
  assign T3796 = T3801 | T6907;
  assign T6907 = {T6909, T3797};
  assign T3797 = T6908 & T3798;
  assign T3798 = 10'h100;
  assign T6908 = T3799 ? 10'h3ff : 10'h0;
  assign T3799 = T3800;
  assign T3800 = 1'h1;
  assign T6909 = T6910 ? 7'h7f : 7'h0;
  assign T6910 = T3797[4'h9];
  assign T3801 = T3723 & T6911;
  assign T6911 = {T6912, T3802};
  assign T3802 = ~ T3798;
  assign T6912 = T6913 ? 7'h7f : 7'h0;
  assign T6913 = T3802[4'h9];
  assign T3803 = T3740 & T3804;
  assign T3804 = 4'h7 == T3739;
  assign T3805 = T3810 | T6914;
  assign T6914 = {T6916, T3806};
  assign T3806 = T6915 & T3807;
  assign T3807 = 9'h80;
  assign T6915 = T3808 ? 9'h1ff : 9'h0;
  assign T3808 = T3809;
  assign T3809 = 1'h1;
  assign T6916 = T6917 ? 8'hff : 8'h0;
  assign T6917 = T3806[4'h8];
  assign T3810 = T3722 & T6918;
  assign T6918 = {T6919, T3811};
  assign T3811 = ~ T3807;
  assign T6919 = T6920 ? 8'hff : 8'h0;
  assign T6920 = T3811[4'h8];
  assign T3812 = T3740 & T3813;
  assign T3813 = 4'h8 == T3739;
  assign T3814 = T3819 | T6921;
  assign T6921 = {T6923, T3815};
  assign T3815 = T6922 & T3816;
  assign T3816 = 8'h40;
  assign T6922 = T3817 ? 8'hff : 8'h0;
  assign T3817 = T3818;
  assign T3818 = 1'h1;
  assign T6923 = T6924 ? 9'h1ff : 9'h0;
  assign T6924 = T3815[3'h7];
  assign T3819 = T3721 & T6925;
  assign T6925 = {T6926, T3820};
  assign T3820 = ~ T3816;
  assign T6926 = T6927 ? 9'h1ff : 9'h0;
  assign T6927 = T3820[3'h7];
  assign T3821 = T3740 & T3822;
  assign T3822 = 4'h9 == T3739;
  assign T3823 = T3828 | T6928;
  assign T6928 = {T6930, T3824};
  assign T3824 = T6929 & T3825;
  assign T3825 = 7'h20;
  assign T6929 = T3826 ? 7'h7f : 7'h0;
  assign T3826 = T3827;
  assign T3827 = 1'h1;
  assign T6930 = T6931 ? 10'h3ff : 10'h0;
  assign T6931 = T3824[3'h6];
  assign T3828 = T3720 & T6932;
  assign T6932 = {T6933, T3829};
  assign T3829 = ~ T3825;
  assign T6933 = T6934 ? 10'h3ff : 10'h0;
  assign T6934 = T3829[3'h6];
  assign T3830 = T3740 & T3831;
  assign T3831 = 4'ha == T3739;
  assign T3832 = T3837 | T6935;
  assign T6935 = {T6937, T3833};
  assign T3833 = T6936 & T3834;
  assign T3834 = 6'h10;
  assign T6936 = T3835 ? 6'h3f : 6'h0;
  assign T3835 = T3836;
  assign T3836 = 1'h1;
  assign T6937 = T6938 ? 11'h7ff : 11'h0;
  assign T6938 = T3833[3'h5];
  assign T3837 = T3719 & T6939;
  assign T6939 = {T6940, T3838};
  assign T3838 = ~ T3834;
  assign T6940 = T6941 ? 11'h7ff : 11'h0;
  assign T6941 = T3838[3'h5];
  assign T3839 = T3740 & T3840;
  assign T3840 = 4'hb == T3739;
  assign T3841 = T3846 | T6942;
  assign T6942 = {T6944, T3842};
  assign T3842 = T6943 & T3843;
  assign T3843 = 5'h8;
  assign T6943 = T3844 ? 5'h1f : 5'h0;
  assign T3844 = T3845;
  assign T3845 = 1'h1;
  assign T6944 = T6945 ? 12'hfff : 12'h0;
  assign T6945 = T3842[3'h4];
  assign T3846 = T3718 & T6946;
  assign T6946 = {T6947, T3847};
  assign T3847 = ~ T3843;
  assign T6947 = T6948 ? 12'hfff : 12'h0;
  assign T6948 = T3847[3'h4];
  assign T3848 = T3740 & T3849;
  assign T3849 = 4'hc == T3739;
  assign T3850 = T3855 | T6949;
  assign T6949 = {T6951, T3851};
  assign T3851 = T6950 & T3852;
  assign T3852 = 4'h4;
  assign T6950 = T3853 ? 4'hf : 4'h0;
  assign T3853 = T3854;
  assign T3854 = 1'h1;
  assign T6951 = T6952 ? 13'h1fff : 13'h0;
  assign T6952 = T3851[2'h3];
  assign T3855 = T3717 & T6953;
  assign T6953 = {T6954, T3856};
  assign T3856 = ~ T3852;
  assign T6954 = T6955 ? 13'h1fff : 13'h0;
  assign T6955 = T3856[2'h3];
  assign T3857 = T3740 & T3858;
  assign T3858 = 4'hd == T3739;
  assign T3859 = T3864 | T6956;
  assign T6956 = {T6958, T3860};
  assign T3860 = T6957 & T3861;
  assign T3861 = 3'h2;
  assign T6957 = T3862 ? 3'h7 : 3'h0;
  assign T3862 = T3863;
  assign T3863 = 1'h1;
  assign T6958 = T6959 ? 14'h3fff : 14'h0;
  assign T6959 = T3860[2'h2];
  assign T3864 = T3716 & T6960;
  assign T6960 = {T6961, T3865};
  assign T3865 = ~ T3861;
  assign T6961 = T6962 ? 14'h3fff : 14'h0;
  assign T6962 = T3865[2'h2];
  assign T3866 = T3740 & T3867;
  assign T3867 = 4'he == T3739;
  assign T3868 = T3873 | T6963;
  assign T6963 = {T6965, T3869};
  assign T3869 = T6964 & T3870;
  assign T3870 = 2'h1;
  assign T6964 = T3871 ? 2'h3 : 2'h0;
  assign T3871 = T3872;
  assign T3872 = 1'h1;
  assign T6965 = T6966 ? 15'h7fff : 15'h0;
  assign T6966 = T3869[1'h1];
  assign T3873 = T3715 & T6967;
  assign T6967 = {T6968, T3874};
  assign T3874 = ~ T3870;
  assign T6968 = T6969 ? 15'h7fff : 15'h0;
  assign T6969 = T3874[1'h1];
  assign T3875 = T3740 & T3876;
  assign T3876 = 4'hf == T3739;
  assign io_V_wire_en_16 = V_wire_en_16;
  assign V_wire_en_16 = T6970;
  assign T6970 = T3877[4'hf:1'h0];
  assign T3877 = T4038 ? T4031 : T3878;
  assign T3878 = T4029 ? T4022 : T3879;
  assign T3879 = T4020 ? T4013 : T3880;
  assign T3880 = T4011 ? T4004 : T3881;
  assign T3881 = T4002 ? T3995 : T3882;
  assign T3882 = T3993 ? T3986 : T3883;
  assign T3883 = T3984 ? T3977 : T3884;
  assign T3884 = T3975 ? T3968 : T3885;
  assign T3885 = T3966 ? T3959 : T3886;
  assign T3886 = T3957 ? T3950 : T3887;
  assign T3887 = T3948 ? T3941 : T3888;
  assign T3888 = T3939 ? T3932 : T3889;
  assign T3889 = T3930 ? T3923 : T3890;
  assign T3890 = T3921 ? T3914 : T3891;
  assign T3891 = T3912 ? T3905 : T3892;
  assign T3892 = T3900 ? T3893 : 17'h0;
  assign T3893 = T3898 | T3894;
  assign T3894 = T6971 & T3895;
  assign T3895 = 17'h8000;
  assign T6971 = T3896 ? 17'h1ffff : 17'h0;
  assign T3896 = T3897;
  assign T3897 = 1'h1;
  assign T3898 = 17'h0 & T3899;
  assign T3899 = ~ T3895;
  assign T3900 = T3903 & T3901;
  assign T3901 = 4'h0 == T3902;
  assign T3902 = LogicBlockModule_16_io_config_V_out[2'h3:1'h0];
  assign T3903 = T3904;
  assign T3904 = LogicBlockModule_16_io_config_V_out[3'h4];
  assign T3905 = T3910 | T6972;
  assign T6972 = {T6974, T3906};
  assign T3906 = T6973 & T3907;
  assign T3907 = 16'h4000;
  assign T6973 = T3908 ? 16'hffff : 16'h0;
  assign T3908 = T3909;
  assign T3909 = 1'h1;
  assign T6974 = T3906[4'hf];
  assign T3910 = T3892 & T6975;
  assign T6975 = {T6976, T3911};
  assign T3911 = ~ T3907;
  assign T6976 = T3911[4'hf];
  assign T3912 = T3903 & T3913;
  assign T3913 = 4'h1 == T3902;
  assign T3914 = T3919 | T6977;
  assign T6977 = {T6979, T3915};
  assign T3915 = T6978 & T3916;
  assign T3916 = 15'h2000;
  assign T6978 = T3917 ? 15'h7fff : 15'h0;
  assign T3917 = T3918;
  assign T3918 = 1'h1;
  assign T6979 = T6980 ? 2'h3 : 2'h0;
  assign T6980 = T3915[4'he];
  assign T3919 = T3891 & T6981;
  assign T6981 = {T6982, T3920};
  assign T3920 = ~ T3916;
  assign T6982 = T6983 ? 2'h3 : 2'h0;
  assign T6983 = T3920[4'he];
  assign T3921 = T3903 & T3922;
  assign T3922 = 4'h2 == T3902;
  assign T3923 = T3928 | T6984;
  assign T6984 = {T6986, T3924};
  assign T3924 = T6985 & T3925;
  assign T3925 = 14'h1000;
  assign T6985 = T3926 ? 14'h3fff : 14'h0;
  assign T3926 = T3927;
  assign T3927 = 1'h1;
  assign T6986 = T6987 ? 3'h7 : 3'h0;
  assign T6987 = T3924[4'hd];
  assign T3928 = T3890 & T6988;
  assign T6988 = {T6989, T3929};
  assign T3929 = ~ T3925;
  assign T6989 = T6990 ? 3'h7 : 3'h0;
  assign T6990 = T3929[4'hd];
  assign T3930 = T3903 & T3931;
  assign T3931 = 4'h3 == T3902;
  assign T3932 = T3937 | T6991;
  assign T6991 = {T6993, T3933};
  assign T3933 = T6992 & T3934;
  assign T3934 = 13'h800;
  assign T6992 = T3935 ? 13'h1fff : 13'h0;
  assign T3935 = T3936;
  assign T3936 = 1'h1;
  assign T6993 = T6994 ? 4'hf : 4'h0;
  assign T6994 = T3933[4'hc];
  assign T3937 = T3889 & T6995;
  assign T6995 = {T6996, T3938};
  assign T3938 = ~ T3934;
  assign T6996 = T6997 ? 4'hf : 4'h0;
  assign T6997 = T3938[4'hc];
  assign T3939 = T3903 & T3940;
  assign T3940 = 4'h4 == T3902;
  assign T3941 = T3946 | T6998;
  assign T6998 = {T7000, T3942};
  assign T3942 = T6999 & T3943;
  assign T3943 = 12'h400;
  assign T6999 = T3944 ? 12'hfff : 12'h0;
  assign T3944 = T3945;
  assign T3945 = 1'h1;
  assign T7000 = T7001 ? 5'h1f : 5'h0;
  assign T7001 = T3942[4'hb];
  assign T3946 = T3888 & T7002;
  assign T7002 = {T7003, T3947};
  assign T3947 = ~ T3943;
  assign T7003 = T7004 ? 5'h1f : 5'h0;
  assign T7004 = T3947[4'hb];
  assign T3948 = T3903 & T3949;
  assign T3949 = 4'h5 == T3902;
  assign T3950 = T3955 | T7005;
  assign T7005 = {T7007, T3951};
  assign T3951 = T7006 & T3952;
  assign T3952 = 11'h200;
  assign T7006 = T3953 ? 11'h7ff : 11'h0;
  assign T3953 = T3954;
  assign T3954 = 1'h1;
  assign T7007 = T7008 ? 6'h3f : 6'h0;
  assign T7008 = T3951[4'ha];
  assign T3955 = T3887 & T7009;
  assign T7009 = {T7010, T3956};
  assign T3956 = ~ T3952;
  assign T7010 = T7011 ? 6'h3f : 6'h0;
  assign T7011 = T3956[4'ha];
  assign T3957 = T3903 & T3958;
  assign T3958 = 4'h6 == T3902;
  assign T3959 = T3964 | T7012;
  assign T7012 = {T7014, T3960};
  assign T3960 = T7013 & T3961;
  assign T3961 = 10'h100;
  assign T7013 = T3962 ? 10'h3ff : 10'h0;
  assign T3962 = T3963;
  assign T3963 = 1'h1;
  assign T7014 = T7015 ? 7'h7f : 7'h0;
  assign T7015 = T3960[4'h9];
  assign T3964 = T3886 & T7016;
  assign T7016 = {T7017, T3965};
  assign T3965 = ~ T3961;
  assign T7017 = T7018 ? 7'h7f : 7'h0;
  assign T7018 = T3965[4'h9];
  assign T3966 = T3903 & T3967;
  assign T3967 = 4'h7 == T3902;
  assign T3968 = T3973 | T7019;
  assign T7019 = {T7021, T3969};
  assign T3969 = T7020 & T3970;
  assign T3970 = 9'h80;
  assign T7020 = T3971 ? 9'h1ff : 9'h0;
  assign T3971 = T3972;
  assign T3972 = 1'h1;
  assign T7021 = T7022 ? 8'hff : 8'h0;
  assign T7022 = T3969[4'h8];
  assign T3973 = T3885 & T7023;
  assign T7023 = {T7024, T3974};
  assign T3974 = ~ T3970;
  assign T7024 = T7025 ? 8'hff : 8'h0;
  assign T7025 = T3974[4'h8];
  assign T3975 = T3903 & T3976;
  assign T3976 = 4'h8 == T3902;
  assign T3977 = T3982 | T7026;
  assign T7026 = {T7028, T3978};
  assign T3978 = T7027 & T3979;
  assign T3979 = 8'h40;
  assign T7027 = T3980 ? 8'hff : 8'h0;
  assign T3980 = T3981;
  assign T3981 = 1'h1;
  assign T7028 = T7029 ? 9'h1ff : 9'h0;
  assign T7029 = T3978[3'h7];
  assign T3982 = T3884 & T7030;
  assign T7030 = {T7031, T3983};
  assign T3983 = ~ T3979;
  assign T7031 = T7032 ? 9'h1ff : 9'h0;
  assign T7032 = T3983[3'h7];
  assign T3984 = T3903 & T3985;
  assign T3985 = 4'h9 == T3902;
  assign T3986 = T3991 | T7033;
  assign T7033 = {T7035, T3987};
  assign T3987 = T7034 & T3988;
  assign T3988 = 7'h20;
  assign T7034 = T3989 ? 7'h7f : 7'h0;
  assign T3989 = T3990;
  assign T3990 = 1'h1;
  assign T7035 = T7036 ? 10'h3ff : 10'h0;
  assign T7036 = T3987[3'h6];
  assign T3991 = T3883 & T7037;
  assign T7037 = {T7038, T3992};
  assign T3992 = ~ T3988;
  assign T7038 = T7039 ? 10'h3ff : 10'h0;
  assign T7039 = T3992[3'h6];
  assign T3993 = T3903 & T3994;
  assign T3994 = 4'ha == T3902;
  assign T3995 = T4000 | T7040;
  assign T7040 = {T7042, T3996};
  assign T3996 = T7041 & T3997;
  assign T3997 = 6'h10;
  assign T7041 = T3998 ? 6'h3f : 6'h0;
  assign T3998 = T3999;
  assign T3999 = 1'h1;
  assign T7042 = T7043 ? 11'h7ff : 11'h0;
  assign T7043 = T3996[3'h5];
  assign T4000 = T3882 & T7044;
  assign T7044 = {T7045, T4001};
  assign T4001 = ~ T3997;
  assign T7045 = T7046 ? 11'h7ff : 11'h0;
  assign T7046 = T4001[3'h5];
  assign T4002 = T3903 & T4003;
  assign T4003 = 4'hb == T3902;
  assign T4004 = T4009 | T7047;
  assign T7047 = {T7049, T4005};
  assign T4005 = T7048 & T4006;
  assign T4006 = 5'h8;
  assign T7048 = T4007 ? 5'h1f : 5'h0;
  assign T4007 = T4008;
  assign T4008 = 1'h1;
  assign T7049 = T7050 ? 12'hfff : 12'h0;
  assign T7050 = T4005[3'h4];
  assign T4009 = T3881 & T7051;
  assign T7051 = {T7052, T4010};
  assign T4010 = ~ T4006;
  assign T7052 = T7053 ? 12'hfff : 12'h0;
  assign T7053 = T4010[3'h4];
  assign T4011 = T3903 & T4012;
  assign T4012 = 4'hc == T3902;
  assign T4013 = T4018 | T7054;
  assign T7054 = {T7056, T4014};
  assign T4014 = T7055 & T4015;
  assign T4015 = 4'h4;
  assign T7055 = T4016 ? 4'hf : 4'h0;
  assign T4016 = T4017;
  assign T4017 = 1'h1;
  assign T7056 = T7057 ? 13'h1fff : 13'h0;
  assign T7057 = T4014[2'h3];
  assign T4018 = T3880 & T7058;
  assign T7058 = {T7059, T4019};
  assign T4019 = ~ T4015;
  assign T7059 = T7060 ? 13'h1fff : 13'h0;
  assign T7060 = T4019[2'h3];
  assign T4020 = T3903 & T4021;
  assign T4021 = 4'hd == T3902;
  assign T4022 = T4027 | T7061;
  assign T7061 = {T7063, T4023};
  assign T4023 = T7062 & T4024;
  assign T4024 = 3'h2;
  assign T7062 = T4025 ? 3'h7 : 3'h0;
  assign T4025 = T4026;
  assign T4026 = 1'h1;
  assign T7063 = T7064 ? 14'h3fff : 14'h0;
  assign T7064 = T4023[2'h2];
  assign T4027 = T3879 & T7065;
  assign T7065 = {T7066, T4028};
  assign T4028 = ~ T4024;
  assign T7066 = T7067 ? 14'h3fff : 14'h0;
  assign T7067 = T4028[2'h2];
  assign T4029 = T3903 & T4030;
  assign T4030 = 4'he == T3902;
  assign T4031 = T4036 | T7068;
  assign T7068 = {T7070, T4032};
  assign T4032 = T7069 & T4033;
  assign T4033 = 2'h1;
  assign T7069 = T4034 ? 2'h3 : 2'h0;
  assign T4034 = T4035;
  assign T4035 = 1'h1;
  assign T7070 = T7071 ? 15'h7fff : 15'h0;
  assign T7071 = T4032[1'h1];
  assign T4036 = T3878 & T7072;
  assign T7072 = {T7073, T4037};
  assign T4037 = ~ T4033;
  assign T7073 = T7074 ? 15'h7fff : 15'h0;
  assign T7074 = T4037[1'h1];
  assign T4038 = T3903 & T4039;
  assign T4039 = 4'hf == T3902;
  assign io_V_wire_en_17 = V_wire_en_17;
  assign V_wire_en_17 = T7075;
  assign T7075 = T4040[4'hf:1'h0];
  assign T4040 = T4201 ? T4194 : T4041;
  assign T4041 = T4192 ? T4185 : T4042;
  assign T4042 = T4183 ? T4176 : T4043;
  assign T4043 = T4174 ? T4167 : T4044;
  assign T4044 = T4165 ? T4158 : T4045;
  assign T4045 = T4156 ? T4149 : T4046;
  assign T4046 = T4147 ? T4140 : T4047;
  assign T4047 = T4138 ? T4131 : T4048;
  assign T4048 = T4129 ? T4122 : T4049;
  assign T4049 = T4120 ? T4113 : T4050;
  assign T4050 = T4111 ? T4104 : T4051;
  assign T4051 = T4102 ? T4095 : T4052;
  assign T4052 = T4093 ? T4086 : T4053;
  assign T4053 = T4084 ? T4077 : T4054;
  assign T4054 = T4075 ? T4068 : T4055;
  assign T4055 = T4063 ? T4056 : 17'h0;
  assign T4056 = T4061 | T4057;
  assign T4057 = T7076 & T4058;
  assign T4058 = 17'h8000;
  assign T7076 = T4059 ? 17'h1ffff : 17'h0;
  assign T4059 = T4060;
  assign T4060 = 1'h1;
  assign T4061 = 17'h0 & T4062;
  assign T4062 = ~ T4058;
  assign T4063 = T4066 & T4064;
  assign T4064 = 4'h0 == T4065;
  assign T4065 = LogicBlockModule_17_io_config_V_out[2'h3:1'h0];
  assign T4066 = T4067;
  assign T4067 = LogicBlockModule_17_io_config_V_out[3'h4];
  assign T4068 = T4073 | T7077;
  assign T7077 = {T7079, T4069};
  assign T4069 = T7078 & T4070;
  assign T4070 = 16'h4000;
  assign T7078 = T4071 ? 16'hffff : 16'h0;
  assign T4071 = T4072;
  assign T4072 = 1'h1;
  assign T7079 = T4069[4'hf];
  assign T4073 = T4055 & T7080;
  assign T7080 = {T7081, T4074};
  assign T4074 = ~ T4070;
  assign T7081 = T4074[4'hf];
  assign T4075 = T4066 & T4076;
  assign T4076 = 4'h1 == T4065;
  assign T4077 = T4082 | T7082;
  assign T7082 = {T7084, T4078};
  assign T4078 = T7083 & T4079;
  assign T4079 = 15'h2000;
  assign T7083 = T4080 ? 15'h7fff : 15'h0;
  assign T4080 = T4081;
  assign T4081 = 1'h1;
  assign T7084 = T7085 ? 2'h3 : 2'h0;
  assign T7085 = T4078[4'he];
  assign T4082 = T4054 & T7086;
  assign T7086 = {T7087, T4083};
  assign T4083 = ~ T4079;
  assign T7087 = T7088 ? 2'h3 : 2'h0;
  assign T7088 = T4083[4'he];
  assign T4084 = T4066 & T4085;
  assign T4085 = 4'h2 == T4065;
  assign T4086 = T4091 | T7089;
  assign T7089 = {T7091, T4087};
  assign T4087 = T7090 & T4088;
  assign T4088 = 14'h1000;
  assign T7090 = T4089 ? 14'h3fff : 14'h0;
  assign T4089 = T4090;
  assign T4090 = 1'h1;
  assign T7091 = T7092 ? 3'h7 : 3'h0;
  assign T7092 = T4087[4'hd];
  assign T4091 = T4053 & T7093;
  assign T7093 = {T7094, T4092};
  assign T4092 = ~ T4088;
  assign T7094 = T7095 ? 3'h7 : 3'h0;
  assign T7095 = T4092[4'hd];
  assign T4093 = T4066 & T4094;
  assign T4094 = 4'h3 == T4065;
  assign T4095 = T4100 | T7096;
  assign T7096 = {T7098, T4096};
  assign T4096 = T7097 & T4097;
  assign T4097 = 13'h800;
  assign T7097 = T4098 ? 13'h1fff : 13'h0;
  assign T4098 = T4099;
  assign T4099 = 1'h1;
  assign T7098 = T7099 ? 4'hf : 4'h0;
  assign T7099 = T4096[4'hc];
  assign T4100 = T4052 & T7100;
  assign T7100 = {T7101, T4101};
  assign T4101 = ~ T4097;
  assign T7101 = T7102 ? 4'hf : 4'h0;
  assign T7102 = T4101[4'hc];
  assign T4102 = T4066 & T4103;
  assign T4103 = 4'h4 == T4065;
  assign T4104 = T4109 | T7103;
  assign T7103 = {T7105, T4105};
  assign T4105 = T7104 & T4106;
  assign T4106 = 12'h400;
  assign T7104 = T4107 ? 12'hfff : 12'h0;
  assign T4107 = T4108;
  assign T4108 = 1'h1;
  assign T7105 = T7106 ? 5'h1f : 5'h0;
  assign T7106 = T4105[4'hb];
  assign T4109 = T4051 & T7107;
  assign T7107 = {T7108, T4110};
  assign T4110 = ~ T4106;
  assign T7108 = T7109 ? 5'h1f : 5'h0;
  assign T7109 = T4110[4'hb];
  assign T4111 = T4066 & T4112;
  assign T4112 = 4'h5 == T4065;
  assign T4113 = T4118 | T7110;
  assign T7110 = {T7112, T4114};
  assign T4114 = T7111 & T4115;
  assign T4115 = 11'h200;
  assign T7111 = T4116 ? 11'h7ff : 11'h0;
  assign T4116 = T4117;
  assign T4117 = 1'h1;
  assign T7112 = T7113 ? 6'h3f : 6'h0;
  assign T7113 = T4114[4'ha];
  assign T4118 = T4050 & T7114;
  assign T7114 = {T7115, T4119};
  assign T4119 = ~ T4115;
  assign T7115 = T7116 ? 6'h3f : 6'h0;
  assign T7116 = T4119[4'ha];
  assign T4120 = T4066 & T4121;
  assign T4121 = 4'h6 == T4065;
  assign T4122 = T4127 | T7117;
  assign T7117 = {T7119, T4123};
  assign T4123 = T7118 & T4124;
  assign T4124 = 10'h100;
  assign T7118 = T4125 ? 10'h3ff : 10'h0;
  assign T4125 = T4126;
  assign T4126 = 1'h1;
  assign T7119 = T7120 ? 7'h7f : 7'h0;
  assign T7120 = T4123[4'h9];
  assign T4127 = T4049 & T7121;
  assign T7121 = {T7122, T4128};
  assign T4128 = ~ T4124;
  assign T7122 = T7123 ? 7'h7f : 7'h0;
  assign T7123 = T4128[4'h9];
  assign T4129 = T4066 & T4130;
  assign T4130 = 4'h7 == T4065;
  assign T4131 = T4136 | T7124;
  assign T7124 = {T7126, T4132};
  assign T4132 = T7125 & T4133;
  assign T4133 = 9'h80;
  assign T7125 = T4134 ? 9'h1ff : 9'h0;
  assign T4134 = T4135;
  assign T4135 = 1'h1;
  assign T7126 = T7127 ? 8'hff : 8'h0;
  assign T7127 = T4132[4'h8];
  assign T4136 = T4048 & T7128;
  assign T7128 = {T7129, T4137};
  assign T4137 = ~ T4133;
  assign T7129 = T7130 ? 8'hff : 8'h0;
  assign T7130 = T4137[4'h8];
  assign T4138 = T4066 & T4139;
  assign T4139 = 4'h8 == T4065;
  assign T4140 = T4145 | T7131;
  assign T7131 = {T7133, T4141};
  assign T4141 = T7132 & T4142;
  assign T4142 = 8'h40;
  assign T7132 = T4143 ? 8'hff : 8'h0;
  assign T4143 = T4144;
  assign T4144 = 1'h1;
  assign T7133 = T7134 ? 9'h1ff : 9'h0;
  assign T7134 = T4141[3'h7];
  assign T4145 = T4047 & T7135;
  assign T7135 = {T7136, T4146};
  assign T4146 = ~ T4142;
  assign T7136 = T7137 ? 9'h1ff : 9'h0;
  assign T7137 = T4146[3'h7];
  assign T4147 = T4066 & T4148;
  assign T4148 = 4'h9 == T4065;
  assign T4149 = T4154 | T7138;
  assign T7138 = {T7140, T4150};
  assign T4150 = T7139 & T4151;
  assign T4151 = 7'h20;
  assign T7139 = T4152 ? 7'h7f : 7'h0;
  assign T4152 = T4153;
  assign T4153 = 1'h1;
  assign T7140 = T7141 ? 10'h3ff : 10'h0;
  assign T7141 = T4150[3'h6];
  assign T4154 = T4046 & T7142;
  assign T7142 = {T7143, T4155};
  assign T4155 = ~ T4151;
  assign T7143 = T7144 ? 10'h3ff : 10'h0;
  assign T7144 = T4155[3'h6];
  assign T4156 = T4066 & T4157;
  assign T4157 = 4'ha == T4065;
  assign T4158 = T4163 | T7145;
  assign T7145 = {T7147, T4159};
  assign T4159 = T7146 & T4160;
  assign T4160 = 6'h10;
  assign T7146 = T4161 ? 6'h3f : 6'h0;
  assign T4161 = T4162;
  assign T4162 = 1'h1;
  assign T7147 = T7148 ? 11'h7ff : 11'h0;
  assign T7148 = T4159[3'h5];
  assign T4163 = T4045 & T7149;
  assign T7149 = {T7150, T4164};
  assign T4164 = ~ T4160;
  assign T7150 = T7151 ? 11'h7ff : 11'h0;
  assign T7151 = T4164[3'h5];
  assign T4165 = T4066 & T4166;
  assign T4166 = 4'hb == T4065;
  assign T4167 = T4172 | T7152;
  assign T7152 = {T7154, T4168};
  assign T4168 = T7153 & T4169;
  assign T4169 = 5'h8;
  assign T7153 = T4170 ? 5'h1f : 5'h0;
  assign T4170 = T4171;
  assign T4171 = 1'h1;
  assign T7154 = T7155 ? 12'hfff : 12'h0;
  assign T7155 = T4168[3'h4];
  assign T4172 = T4044 & T7156;
  assign T7156 = {T7157, T4173};
  assign T4173 = ~ T4169;
  assign T7157 = T7158 ? 12'hfff : 12'h0;
  assign T7158 = T4173[3'h4];
  assign T4174 = T4066 & T4175;
  assign T4175 = 4'hc == T4065;
  assign T4176 = T4181 | T7159;
  assign T7159 = {T7161, T4177};
  assign T4177 = T7160 & T4178;
  assign T4178 = 4'h4;
  assign T7160 = T4179 ? 4'hf : 4'h0;
  assign T4179 = T4180;
  assign T4180 = 1'h1;
  assign T7161 = T7162 ? 13'h1fff : 13'h0;
  assign T7162 = T4177[2'h3];
  assign T4181 = T4043 & T7163;
  assign T7163 = {T7164, T4182};
  assign T4182 = ~ T4178;
  assign T7164 = T7165 ? 13'h1fff : 13'h0;
  assign T7165 = T4182[2'h3];
  assign T4183 = T4066 & T4184;
  assign T4184 = 4'hd == T4065;
  assign T4185 = T4190 | T7166;
  assign T7166 = {T7168, T4186};
  assign T4186 = T7167 & T4187;
  assign T4187 = 3'h2;
  assign T7167 = T4188 ? 3'h7 : 3'h0;
  assign T4188 = T4189;
  assign T4189 = 1'h1;
  assign T7168 = T7169 ? 14'h3fff : 14'h0;
  assign T7169 = T4186[2'h2];
  assign T4190 = T4042 & T7170;
  assign T7170 = {T7171, T4191};
  assign T4191 = ~ T4187;
  assign T7171 = T7172 ? 14'h3fff : 14'h0;
  assign T7172 = T4191[2'h2];
  assign T4192 = T4066 & T4193;
  assign T4193 = 4'he == T4065;
  assign T4194 = T4199 | T7173;
  assign T7173 = {T7175, T4195};
  assign T4195 = T7174 & T4196;
  assign T4196 = 2'h1;
  assign T7174 = T4197 ? 2'h3 : 2'h0;
  assign T4197 = T4198;
  assign T4198 = 1'h1;
  assign T7175 = T7176 ? 15'h7fff : 15'h0;
  assign T7176 = T4195[1'h1];
  assign T4199 = T4041 & T7177;
  assign T7177 = {T7178, T4200};
  assign T4200 = ~ T4196;
  assign T7178 = T7179 ? 15'h7fff : 15'h0;
  assign T7179 = T4200[1'h1];
  assign T4201 = T4066 & T4202;
  assign T4202 = 4'hf == T4065;
  assign io_V_wire_en_18 = V_wire_en_18;
  assign V_wire_en_18 = T7180;
  assign T7180 = T4203[4'hf:1'h0];
  assign T4203 = T4364 ? T4357 : T4204;
  assign T4204 = T4355 ? T4348 : T4205;
  assign T4205 = T4346 ? T4339 : T4206;
  assign T4206 = T4337 ? T4330 : T4207;
  assign T4207 = T4328 ? T4321 : T4208;
  assign T4208 = T4319 ? T4312 : T4209;
  assign T4209 = T4310 ? T4303 : T4210;
  assign T4210 = T4301 ? T4294 : T4211;
  assign T4211 = T4292 ? T4285 : T4212;
  assign T4212 = T4283 ? T4276 : T4213;
  assign T4213 = T4274 ? T4267 : T4214;
  assign T4214 = T4265 ? T4258 : T4215;
  assign T4215 = T4256 ? T4249 : T4216;
  assign T4216 = T4247 ? T4240 : T4217;
  assign T4217 = T4238 ? T4231 : T4218;
  assign T4218 = T4226 ? T4219 : 17'h0;
  assign T4219 = T4224 | T4220;
  assign T4220 = T7181 & T4221;
  assign T4221 = 17'h8000;
  assign T7181 = T4222 ? 17'h1ffff : 17'h0;
  assign T4222 = T4223;
  assign T4223 = 1'h1;
  assign T4224 = 17'h0 & T4225;
  assign T4225 = ~ T4221;
  assign T4226 = T4229 & T4227;
  assign T4227 = 4'h0 == T4228;
  assign T4228 = LogicBlockModule_18_io_config_V_out[2'h3:1'h0];
  assign T4229 = T4230;
  assign T4230 = LogicBlockModule_18_io_config_V_out[3'h4];
  assign T4231 = T4236 | T7182;
  assign T7182 = {T7184, T4232};
  assign T4232 = T7183 & T4233;
  assign T4233 = 16'h4000;
  assign T7183 = T4234 ? 16'hffff : 16'h0;
  assign T4234 = T4235;
  assign T4235 = 1'h1;
  assign T7184 = T4232[4'hf];
  assign T4236 = T4218 & T7185;
  assign T7185 = {T7186, T4237};
  assign T4237 = ~ T4233;
  assign T7186 = T4237[4'hf];
  assign T4238 = T4229 & T4239;
  assign T4239 = 4'h1 == T4228;
  assign T4240 = T4245 | T7187;
  assign T7187 = {T7189, T4241};
  assign T4241 = T7188 & T4242;
  assign T4242 = 15'h2000;
  assign T7188 = T4243 ? 15'h7fff : 15'h0;
  assign T4243 = T4244;
  assign T4244 = 1'h1;
  assign T7189 = T7190 ? 2'h3 : 2'h0;
  assign T7190 = T4241[4'he];
  assign T4245 = T4217 & T7191;
  assign T7191 = {T7192, T4246};
  assign T4246 = ~ T4242;
  assign T7192 = T7193 ? 2'h3 : 2'h0;
  assign T7193 = T4246[4'he];
  assign T4247 = T4229 & T4248;
  assign T4248 = 4'h2 == T4228;
  assign T4249 = T4254 | T7194;
  assign T7194 = {T7196, T4250};
  assign T4250 = T7195 & T4251;
  assign T4251 = 14'h1000;
  assign T7195 = T4252 ? 14'h3fff : 14'h0;
  assign T4252 = T4253;
  assign T4253 = 1'h1;
  assign T7196 = T7197 ? 3'h7 : 3'h0;
  assign T7197 = T4250[4'hd];
  assign T4254 = T4216 & T7198;
  assign T7198 = {T7199, T4255};
  assign T4255 = ~ T4251;
  assign T7199 = T7200 ? 3'h7 : 3'h0;
  assign T7200 = T4255[4'hd];
  assign T4256 = T4229 & T4257;
  assign T4257 = 4'h3 == T4228;
  assign T4258 = T4263 | T7201;
  assign T7201 = {T7203, T4259};
  assign T4259 = T7202 & T4260;
  assign T4260 = 13'h800;
  assign T7202 = T4261 ? 13'h1fff : 13'h0;
  assign T4261 = T4262;
  assign T4262 = 1'h1;
  assign T7203 = T7204 ? 4'hf : 4'h0;
  assign T7204 = T4259[4'hc];
  assign T4263 = T4215 & T7205;
  assign T7205 = {T7206, T4264};
  assign T4264 = ~ T4260;
  assign T7206 = T7207 ? 4'hf : 4'h0;
  assign T7207 = T4264[4'hc];
  assign T4265 = T4229 & T4266;
  assign T4266 = 4'h4 == T4228;
  assign T4267 = T4272 | T7208;
  assign T7208 = {T7210, T4268};
  assign T4268 = T7209 & T4269;
  assign T4269 = 12'h400;
  assign T7209 = T4270 ? 12'hfff : 12'h0;
  assign T4270 = T4271;
  assign T4271 = 1'h1;
  assign T7210 = T7211 ? 5'h1f : 5'h0;
  assign T7211 = T4268[4'hb];
  assign T4272 = T4214 & T7212;
  assign T7212 = {T7213, T4273};
  assign T4273 = ~ T4269;
  assign T7213 = T7214 ? 5'h1f : 5'h0;
  assign T7214 = T4273[4'hb];
  assign T4274 = T4229 & T4275;
  assign T4275 = 4'h5 == T4228;
  assign T4276 = T4281 | T7215;
  assign T7215 = {T7217, T4277};
  assign T4277 = T7216 & T4278;
  assign T4278 = 11'h200;
  assign T7216 = T4279 ? 11'h7ff : 11'h0;
  assign T4279 = T4280;
  assign T4280 = 1'h1;
  assign T7217 = T7218 ? 6'h3f : 6'h0;
  assign T7218 = T4277[4'ha];
  assign T4281 = T4213 & T7219;
  assign T7219 = {T7220, T4282};
  assign T4282 = ~ T4278;
  assign T7220 = T7221 ? 6'h3f : 6'h0;
  assign T7221 = T4282[4'ha];
  assign T4283 = T4229 & T4284;
  assign T4284 = 4'h6 == T4228;
  assign T4285 = T4290 | T7222;
  assign T7222 = {T7224, T4286};
  assign T4286 = T7223 & T4287;
  assign T4287 = 10'h100;
  assign T7223 = T4288 ? 10'h3ff : 10'h0;
  assign T4288 = T4289;
  assign T4289 = 1'h1;
  assign T7224 = T7225 ? 7'h7f : 7'h0;
  assign T7225 = T4286[4'h9];
  assign T4290 = T4212 & T7226;
  assign T7226 = {T7227, T4291};
  assign T4291 = ~ T4287;
  assign T7227 = T7228 ? 7'h7f : 7'h0;
  assign T7228 = T4291[4'h9];
  assign T4292 = T4229 & T4293;
  assign T4293 = 4'h7 == T4228;
  assign T4294 = T4299 | T7229;
  assign T7229 = {T7231, T4295};
  assign T4295 = T7230 & T4296;
  assign T4296 = 9'h80;
  assign T7230 = T4297 ? 9'h1ff : 9'h0;
  assign T4297 = T4298;
  assign T4298 = 1'h1;
  assign T7231 = T7232 ? 8'hff : 8'h0;
  assign T7232 = T4295[4'h8];
  assign T4299 = T4211 & T7233;
  assign T7233 = {T7234, T4300};
  assign T4300 = ~ T4296;
  assign T7234 = T7235 ? 8'hff : 8'h0;
  assign T7235 = T4300[4'h8];
  assign T4301 = T4229 & T4302;
  assign T4302 = 4'h8 == T4228;
  assign T4303 = T4308 | T7236;
  assign T7236 = {T7238, T4304};
  assign T4304 = T7237 & T4305;
  assign T4305 = 8'h40;
  assign T7237 = T4306 ? 8'hff : 8'h0;
  assign T4306 = T4307;
  assign T4307 = 1'h1;
  assign T7238 = T7239 ? 9'h1ff : 9'h0;
  assign T7239 = T4304[3'h7];
  assign T4308 = T4210 & T7240;
  assign T7240 = {T7241, T4309};
  assign T4309 = ~ T4305;
  assign T7241 = T7242 ? 9'h1ff : 9'h0;
  assign T7242 = T4309[3'h7];
  assign T4310 = T4229 & T4311;
  assign T4311 = 4'h9 == T4228;
  assign T4312 = T4317 | T7243;
  assign T7243 = {T7245, T4313};
  assign T4313 = T7244 & T4314;
  assign T4314 = 7'h20;
  assign T7244 = T4315 ? 7'h7f : 7'h0;
  assign T4315 = T4316;
  assign T4316 = 1'h1;
  assign T7245 = T7246 ? 10'h3ff : 10'h0;
  assign T7246 = T4313[3'h6];
  assign T4317 = T4209 & T7247;
  assign T7247 = {T7248, T4318};
  assign T4318 = ~ T4314;
  assign T7248 = T7249 ? 10'h3ff : 10'h0;
  assign T7249 = T4318[3'h6];
  assign T4319 = T4229 & T4320;
  assign T4320 = 4'ha == T4228;
  assign T4321 = T4326 | T7250;
  assign T7250 = {T7252, T4322};
  assign T4322 = T7251 & T4323;
  assign T4323 = 6'h10;
  assign T7251 = T4324 ? 6'h3f : 6'h0;
  assign T4324 = T4325;
  assign T4325 = 1'h1;
  assign T7252 = T7253 ? 11'h7ff : 11'h0;
  assign T7253 = T4322[3'h5];
  assign T4326 = T4208 & T7254;
  assign T7254 = {T7255, T4327};
  assign T4327 = ~ T4323;
  assign T7255 = T7256 ? 11'h7ff : 11'h0;
  assign T7256 = T4327[3'h5];
  assign T4328 = T4229 & T4329;
  assign T4329 = 4'hb == T4228;
  assign T4330 = T4335 | T7257;
  assign T7257 = {T7259, T4331};
  assign T4331 = T7258 & T4332;
  assign T4332 = 5'h8;
  assign T7258 = T4333 ? 5'h1f : 5'h0;
  assign T4333 = T4334;
  assign T4334 = 1'h1;
  assign T7259 = T7260 ? 12'hfff : 12'h0;
  assign T7260 = T4331[3'h4];
  assign T4335 = T4207 & T7261;
  assign T7261 = {T7262, T4336};
  assign T4336 = ~ T4332;
  assign T7262 = T7263 ? 12'hfff : 12'h0;
  assign T7263 = T4336[3'h4];
  assign T4337 = T4229 & T4338;
  assign T4338 = 4'hc == T4228;
  assign T4339 = T4344 | T7264;
  assign T7264 = {T7266, T4340};
  assign T4340 = T7265 & T4341;
  assign T4341 = 4'h4;
  assign T7265 = T4342 ? 4'hf : 4'h0;
  assign T4342 = T4343;
  assign T4343 = 1'h1;
  assign T7266 = T7267 ? 13'h1fff : 13'h0;
  assign T7267 = T4340[2'h3];
  assign T4344 = T4206 & T7268;
  assign T7268 = {T7269, T4345};
  assign T4345 = ~ T4341;
  assign T7269 = T7270 ? 13'h1fff : 13'h0;
  assign T7270 = T4345[2'h3];
  assign T4346 = T4229 & T4347;
  assign T4347 = 4'hd == T4228;
  assign T4348 = T4353 | T7271;
  assign T7271 = {T7273, T4349};
  assign T4349 = T7272 & T4350;
  assign T4350 = 3'h2;
  assign T7272 = T4351 ? 3'h7 : 3'h0;
  assign T4351 = T4352;
  assign T4352 = 1'h1;
  assign T7273 = T7274 ? 14'h3fff : 14'h0;
  assign T7274 = T4349[2'h2];
  assign T4353 = T4205 & T7275;
  assign T7275 = {T7276, T4354};
  assign T4354 = ~ T4350;
  assign T7276 = T7277 ? 14'h3fff : 14'h0;
  assign T7277 = T4354[2'h2];
  assign T4355 = T4229 & T4356;
  assign T4356 = 4'he == T4228;
  assign T4357 = T4362 | T7278;
  assign T7278 = {T7280, T4358};
  assign T4358 = T7279 & T4359;
  assign T4359 = 2'h1;
  assign T7279 = T4360 ? 2'h3 : 2'h0;
  assign T4360 = T4361;
  assign T4361 = 1'h1;
  assign T7280 = T7281 ? 15'h7fff : 15'h0;
  assign T7281 = T4358[1'h1];
  assign T4362 = T4204 & T7282;
  assign T7282 = {T7283, T4363};
  assign T4363 = ~ T4359;
  assign T7283 = T7284 ? 15'h7fff : 15'h0;
  assign T7284 = T4363[1'h1];
  assign T4364 = T4229 & T4365;
  assign T4365 = 4'hf == T4228;
  assign io_V_wire_en_19 = V_wire_en_19;
  assign V_wire_en_19 = T7285;
  assign T7285 = T4366[4'hf:1'h0];
  assign T4366 = T4527 ? T4520 : T4367;
  assign T4367 = T4518 ? T4511 : T4368;
  assign T4368 = T4509 ? T4502 : T4369;
  assign T4369 = T4500 ? T4493 : T4370;
  assign T4370 = T4491 ? T4484 : T4371;
  assign T4371 = T4482 ? T4475 : T4372;
  assign T4372 = T4473 ? T4466 : T4373;
  assign T4373 = T4464 ? T4457 : T4374;
  assign T4374 = T4455 ? T4448 : T4375;
  assign T4375 = T4446 ? T4439 : T4376;
  assign T4376 = T4437 ? T4430 : T4377;
  assign T4377 = T4428 ? T4421 : T4378;
  assign T4378 = T4419 ? T4412 : T4379;
  assign T4379 = T4410 ? T4403 : T4380;
  assign T4380 = T4401 ? T4394 : T4381;
  assign T4381 = T4389 ? T4382 : 17'h0;
  assign T4382 = T4387 | T4383;
  assign T4383 = T7286 & T4384;
  assign T4384 = 17'h8000;
  assign T7286 = T4385 ? 17'h1ffff : 17'h0;
  assign T4385 = T4386;
  assign T4386 = 1'h1;
  assign T4387 = 17'h0 & T4388;
  assign T4388 = ~ T4384;
  assign T4389 = T4392 & T4390;
  assign T4390 = 4'h0 == T4391;
  assign T4391 = LogicBlockModule_19_io_config_V_out[2'h3:1'h0];
  assign T4392 = T4393;
  assign T4393 = LogicBlockModule_19_io_config_V_out[3'h4];
  assign T4394 = T4399 | T7287;
  assign T7287 = {T7289, T4395};
  assign T4395 = T7288 & T4396;
  assign T4396 = 16'h4000;
  assign T7288 = T4397 ? 16'hffff : 16'h0;
  assign T4397 = T4398;
  assign T4398 = 1'h1;
  assign T7289 = T4395[4'hf];
  assign T4399 = T4381 & T7290;
  assign T7290 = {T7291, T4400};
  assign T4400 = ~ T4396;
  assign T7291 = T4400[4'hf];
  assign T4401 = T4392 & T4402;
  assign T4402 = 4'h1 == T4391;
  assign T4403 = T4408 | T7292;
  assign T7292 = {T7294, T4404};
  assign T4404 = T7293 & T4405;
  assign T4405 = 15'h2000;
  assign T7293 = T4406 ? 15'h7fff : 15'h0;
  assign T4406 = T4407;
  assign T4407 = 1'h1;
  assign T7294 = T7295 ? 2'h3 : 2'h0;
  assign T7295 = T4404[4'he];
  assign T4408 = T4380 & T7296;
  assign T7296 = {T7297, T4409};
  assign T4409 = ~ T4405;
  assign T7297 = T7298 ? 2'h3 : 2'h0;
  assign T7298 = T4409[4'he];
  assign T4410 = T4392 & T4411;
  assign T4411 = 4'h2 == T4391;
  assign T4412 = T4417 | T7299;
  assign T7299 = {T7301, T4413};
  assign T4413 = T7300 & T4414;
  assign T4414 = 14'h1000;
  assign T7300 = T4415 ? 14'h3fff : 14'h0;
  assign T4415 = T4416;
  assign T4416 = 1'h1;
  assign T7301 = T7302 ? 3'h7 : 3'h0;
  assign T7302 = T4413[4'hd];
  assign T4417 = T4379 & T7303;
  assign T7303 = {T7304, T4418};
  assign T4418 = ~ T4414;
  assign T7304 = T7305 ? 3'h7 : 3'h0;
  assign T7305 = T4418[4'hd];
  assign T4419 = T4392 & T4420;
  assign T4420 = 4'h3 == T4391;
  assign T4421 = T4426 | T7306;
  assign T7306 = {T7308, T4422};
  assign T4422 = T7307 & T4423;
  assign T4423 = 13'h800;
  assign T7307 = T4424 ? 13'h1fff : 13'h0;
  assign T4424 = T4425;
  assign T4425 = 1'h1;
  assign T7308 = T7309 ? 4'hf : 4'h0;
  assign T7309 = T4422[4'hc];
  assign T4426 = T4378 & T7310;
  assign T7310 = {T7311, T4427};
  assign T4427 = ~ T4423;
  assign T7311 = T7312 ? 4'hf : 4'h0;
  assign T7312 = T4427[4'hc];
  assign T4428 = T4392 & T4429;
  assign T4429 = 4'h4 == T4391;
  assign T4430 = T4435 | T7313;
  assign T7313 = {T7315, T4431};
  assign T4431 = T7314 & T4432;
  assign T4432 = 12'h400;
  assign T7314 = T4433 ? 12'hfff : 12'h0;
  assign T4433 = T4434;
  assign T4434 = 1'h1;
  assign T7315 = T7316 ? 5'h1f : 5'h0;
  assign T7316 = T4431[4'hb];
  assign T4435 = T4377 & T7317;
  assign T7317 = {T7318, T4436};
  assign T4436 = ~ T4432;
  assign T7318 = T7319 ? 5'h1f : 5'h0;
  assign T7319 = T4436[4'hb];
  assign T4437 = T4392 & T4438;
  assign T4438 = 4'h5 == T4391;
  assign T4439 = T4444 | T7320;
  assign T7320 = {T7322, T4440};
  assign T4440 = T7321 & T4441;
  assign T4441 = 11'h200;
  assign T7321 = T4442 ? 11'h7ff : 11'h0;
  assign T4442 = T4443;
  assign T4443 = 1'h1;
  assign T7322 = T7323 ? 6'h3f : 6'h0;
  assign T7323 = T4440[4'ha];
  assign T4444 = T4376 & T7324;
  assign T7324 = {T7325, T4445};
  assign T4445 = ~ T4441;
  assign T7325 = T7326 ? 6'h3f : 6'h0;
  assign T7326 = T4445[4'ha];
  assign T4446 = T4392 & T4447;
  assign T4447 = 4'h6 == T4391;
  assign T4448 = T4453 | T7327;
  assign T7327 = {T7329, T4449};
  assign T4449 = T7328 & T4450;
  assign T4450 = 10'h100;
  assign T7328 = T4451 ? 10'h3ff : 10'h0;
  assign T4451 = T4452;
  assign T4452 = 1'h1;
  assign T7329 = T7330 ? 7'h7f : 7'h0;
  assign T7330 = T4449[4'h9];
  assign T4453 = T4375 & T7331;
  assign T7331 = {T7332, T4454};
  assign T4454 = ~ T4450;
  assign T7332 = T7333 ? 7'h7f : 7'h0;
  assign T7333 = T4454[4'h9];
  assign T4455 = T4392 & T4456;
  assign T4456 = 4'h7 == T4391;
  assign T4457 = T4462 | T7334;
  assign T7334 = {T7336, T4458};
  assign T4458 = T7335 & T4459;
  assign T4459 = 9'h80;
  assign T7335 = T4460 ? 9'h1ff : 9'h0;
  assign T4460 = T4461;
  assign T4461 = 1'h1;
  assign T7336 = T7337 ? 8'hff : 8'h0;
  assign T7337 = T4458[4'h8];
  assign T4462 = T4374 & T7338;
  assign T7338 = {T7339, T4463};
  assign T4463 = ~ T4459;
  assign T7339 = T7340 ? 8'hff : 8'h0;
  assign T7340 = T4463[4'h8];
  assign T4464 = T4392 & T4465;
  assign T4465 = 4'h8 == T4391;
  assign T4466 = T4471 | T7341;
  assign T7341 = {T7343, T4467};
  assign T4467 = T7342 & T4468;
  assign T4468 = 8'h40;
  assign T7342 = T4469 ? 8'hff : 8'h0;
  assign T4469 = T4470;
  assign T4470 = 1'h1;
  assign T7343 = T7344 ? 9'h1ff : 9'h0;
  assign T7344 = T4467[3'h7];
  assign T4471 = T4373 & T7345;
  assign T7345 = {T7346, T4472};
  assign T4472 = ~ T4468;
  assign T7346 = T7347 ? 9'h1ff : 9'h0;
  assign T7347 = T4472[3'h7];
  assign T4473 = T4392 & T4474;
  assign T4474 = 4'h9 == T4391;
  assign T4475 = T4480 | T7348;
  assign T7348 = {T7350, T4476};
  assign T4476 = T7349 & T4477;
  assign T4477 = 7'h20;
  assign T7349 = T4478 ? 7'h7f : 7'h0;
  assign T4478 = T4479;
  assign T4479 = 1'h1;
  assign T7350 = T7351 ? 10'h3ff : 10'h0;
  assign T7351 = T4476[3'h6];
  assign T4480 = T4372 & T7352;
  assign T7352 = {T7353, T4481};
  assign T4481 = ~ T4477;
  assign T7353 = T7354 ? 10'h3ff : 10'h0;
  assign T7354 = T4481[3'h6];
  assign T4482 = T4392 & T4483;
  assign T4483 = 4'ha == T4391;
  assign T4484 = T4489 | T7355;
  assign T7355 = {T7357, T4485};
  assign T4485 = T7356 & T4486;
  assign T4486 = 6'h10;
  assign T7356 = T4487 ? 6'h3f : 6'h0;
  assign T4487 = T4488;
  assign T4488 = 1'h1;
  assign T7357 = T7358 ? 11'h7ff : 11'h0;
  assign T7358 = T4485[3'h5];
  assign T4489 = T4371 & T7359;
  assign T7359 = {T7360, T4490};
  assign T4490 = ~ T4486;
  assign T7360 = T7361 ? 11'h7ff : 11'h0;
  assign T7361 = T4490[3'h5];
  assign T4491 = T4392 & T4492;
  assign T4492 = 4'hb == T4391;
  assign T4493 = T4498 | T7362;
  assign T7362 = {T7364, T4494};
  assign T4494 = T7363 & T4495;
  assign T4495 = 5'h8;
  assign T7363 = T4496 ? 5'h1f : 5'h0;
  assign T4496 = T4497;
  assign T4497 = 1'h1;
  assign T7364 = T7365 ? 12'hfff : 12'h0;
  assign T7365 = T4494[3'h4];
  assign T4498 = T4370 & T7366;
  assign T7366 = {T7367, T4499};
  assign T4499 = ~ T4495;
  assign T7367 = T7368 ? 12'hfff : 12'h0;
  assign T7368 = T4499[3'h4];
  assign T4500 = T4392 & T4501;
  assign T4501 = 4'hc == T4391;
  assign T4502 = T4507 | T7369;
  assign T7369 = {T7371, T4503};
  assign T4503 = T7370 & T4504;
  assign T4504 = 4'h4;
  assign T7370 = T4505 ? 4'hf : 4'h0;
  assign T4505 = T4506;
  assign T4506 = 1'h1;
  assign T7371 = T7372 ? 13'h1fff : 13'h0;
  assign T7372 = T4503[2'h3];
  assign T4507 = T4369 & T7373;
  assign T7373 = {T7374, T4508};
  assign T4508 = ~ T4504;
  assign T7374 = T7375 ? 13'h1fff : 13'h0;
  assign T7375 = T4508[2'h3];
  assign T4509 = T4392 & T4510;
  assign T4510 = 4'hd == T4391;
  assign T4511 = T4516 | T7376;
  assign T7376 = {T7378, T4512};
  assign T4512 = T7377 & T4513;
  assign T4513 = 3'h2;
  assign T7377 = T4514 ? 3'h7 : 3'h0;
  assign T4514 = T4515;
  assign T4515 = 1'h1;
  assign T7378 = T7379 ? 14'h3fff : 14'h0;
  assign T7379 = T4512[2'h2];
  assign T4516 = T4368 & T7380;
  assign T7380 = {T7381, T4517};
  assign T4517 = ~ T4513;
  assign T7381 = T7382 ? 14'h3fff : 14'h0;
  assign T7382 = T4517[2'h2];
  assign T4518 = T4392 & T4519;
  assign T4519 = 4'he == T4391;
  assign T4520 = T4525 | T7383;
  assign T7383 = {T7385, T4521};
  assign T4521 = T7384 & T4522;
  assign T4522 = 2'h1;
  assign T7384 = T4523 ? 2'h3 : 2'h0;
  assign T4523 = T4524;
  assign T4524 = 1'h1;
  assign T7385 = T7386 ? 15'h7fff : 15'h0;
  assign T7386 = T4521[1'h1];
  assign T4525 = T4367 & T7387;
  assign T7387 = {T7388, T4526};
  assign T4526 = ~ T4522;
  assign T7388 = T7389 ? 15'h7fff : 15'h0;
  assign T7389 = T4526[1'h1];
  assign T4527 = T4392 & T4528;
  assign T4528 = 4'hf == T4391;
  assign io_V_wire_en_20 = V_wire_en_20;
  assign V_wire_en_20 = T7390;
  assign T7390 = T4529[4'hf:1'h0];
  assign T4529 = T4690 ? T4683 : T4530;
  assign T4530 = T4681 ? T4674 : T4531;
  assign T4531 = T4672 ? T4665 : T4532;
  assign T4532 = T4663 ? T4656 : T4533;
  assign T4533 = T4654 ? T4647 : T4534;
  assign T4534 = T4645 ? T4638 : T4535;
  assign T4535 = T4636 ? T4629 : T4536;
  assign T4536 = T4627 ? T4620 : T4537;
  assign T4537 = T4618 ? T4611 : T4538;
  assign T4538 = T4609 ? T4602 : T4539;
  assign T4539 = T4600 ? T4593 : T4540;
  assign T4540 = T4591 ? T4584 : T4541;
  assign T4541 = T4582 ? T4575 : T4542;
  assign T4542 = T4573 ? T4566 : T4543;
  assign T4543 = T4564 ? T4557 : T4544;
  assign T4544 = T4552 ? T4545 : 17'h0;
  assign T4545 = T4550 | T4546;
  assign T4546 = T7391 & T4547;
  assign T4547 = 17'h8000;
  assign T7391 = T4548 ? 17'h1ffff : 17'h0;
  assign T4548 = T4549;
  assign T4549 = 1'h1;
  assign T4550 = 17'h0 & T4551;
  assign T4551 = ~ T4547;
  assign T4552 = T4555 & T4553;
  assign T4553 = 4'h0 == T4554;
  assign T4554 = LogicBlockModule_20_io_config_V_out[2'h3:1'h0];
  assign T4555 = T4556;
  assign T4556 = LogicBlockModule_20_io_config_V_out[3'h4];
  assign T4557 = T4562 | T7392;
  assign T7392 = {T7394, T4558};
  assign T4558 = T7393 & T4559;
  assign T4559 = 16'h4000;
  assign T7393 = T4560 ? 16'hffff : 16'h0;
  assign T4560 = T4561;
  assign T4561 = 1'h1;
  assign T7394 = T4558[4'hf];
  assign T4562 = T4544 & T7395;
  assign T7395 = {T7396, T4563};
  assign T4563 = ~ T4559;
  assign T7396 = T4563[4'hf];
  assign T4564 = T4555 & T4565;
  assign T4565 = 4'h1 == T4554;
  assign T4566 = T4571 | T7397;
  assign T7397 = {T7399, T4567};
  assign T4567 = T7398 & T4568;
  assign T4568 = 15'h2000;
  assign T7398 = T4569 ? 15'h7fff : 15'h0;
  assign T4569 = T4570;
  assign T4570 = 1'h1;
  assign T7399 = T7400 ? 2'h3 : 2'h0;
  assign T7400 = T4567[4'he];
  assign T4571 = T4543 & T7401;
  assign T7401 = {T7402, T4572};
  assign T4572 = ~ T4568;
  assign T7402 = T7403 ? 2'h3 : 2'h0;
  assign T7403 = T4572[4'he];
  assign T4573 = T4555 & T4574;
  assign T4574 = 4'h2 == T4554;
  assign T4575 = T4580 | T7404;
  assign T7404 = {T7406, T4576};
  assign T4576 = T7405 & T4577;
  assign T4577 = 14'h1000;
  assign T7405 = T4578 ? 14'h3fff : 14'h0;
  assign T4578 = T4579;
  assign T4579 = 1'h1;
  assign T7406 = T7407 ? 3'h7 : 3'h0;
  assign T7407 = T4576[4'hd];
  assign T4580 = T4542 & T7408;
  assign T7408 = {T7409, T4581};
  assign T4581 = ~ T4577;
  assign T7409 = T7410 ? 3'h7 : 3'h0;
  assign T7410 = T4581[4'hd];
  assign T4582 = T4555 & T4583;
  assign T4583 = 4'h3 == T4554;
  assign T4584 = T4589 | T7411;
  assign T7411 = {T7413, T4585};
  assign T4585 = T7412 & T4586;
  assign T4586 = 13'h800;
  assign T7412 = T4587 ? 13'h1fff : 13'h0;
  assign T4587 = T4588;
  assign T4588 = 1'h1;
  assign T7413 = T7414 ? 4'hf : 4'h0;
  assign T7414 = T4585[4'hc];
  assign T4589 = T4541 & T7415;
  assign T7415 = {T7416, T4590};
  assign T4590 = ~ T4586;
  assign T7416 = T7417 ? 4'hf : 4'h0;
  assign T7417 = T4590[4'hc];
  assign T4591 = T4555 & T4592;
  assign T4592 = 4'h4 == T4554;
  assign T4593 = T4598 | T7418;
  assign T7418 = {T7420, T4594};
  assign T4594 = T7419 & T4595;
  assign T4595 = 12'h400;
  assign T7419 = T4596 ? 12'hfff : 12'h0;
  assign T4596 = T4597;
  assign T4597 = 1'h1;
  assign T7420 = T7421 ? 5'h1f : 5'h0;
  assign T7421 = T4594[4'hb];
  assign T4598 = T4540 & T7422;
  assign T7422 = {T7423, T4599};
  assign T4599 = ~ T4595;
  assign T7423 = T7424 ? 5'h1f : 5'h0;
  assign T7424 = T4599[4'hb];
  assign T4600 = T4555 & T4601;
  assign T4601 = 4'h5 == T4554;
  assign T4602 = T4607 | T7425;
  assign T7425 = {T7427, T4603};
  assign T4603 = T7426 & T4604;
  assign T4604 = 11'h200;
  assign T7426 = T4605 ? 11'h7ff : 11'h0;
  assign T4605 = T4606;
  assign T4606 = 1'h1;
  assign T7427 = T7428 ? 6'h3f : 6'h0;
  assign T7428 = T4603[4'ha];
  assign T4607 = T4539 & T7429;
  assign T7429 = {T7430, T4608};
  assign T4608 = ~ T4604;
  assign T7430 = T7431 ? 6'h3f : 6'h0;
  assign T7431 = T4608[4'ha];
  assign T4609 = T4555 & T4610;
  assign T4610 = 4'h6 == T4554;
  assign T4611 = T4616 | T7432;
  assign T7432 = {T7434, T4612};
  assign T4612 = T7433 & T4613;
  assign T4613 = 10'h100;
  assign T7433 = T4614 ? 10'h3ff : 10'h0;
  assign T4614 = T4615;
  assign T4615 = 1'h1;
  assign T7434 = T7435 ? 7'h7f : 7'h0;
  assign T7435 = T4612[4'h9];
  assign T4616 = T4538 & T7436;
  assign T7436 = {T7437, T4617};
  assign T4617 = ~ T4613;
  assign T7437 = T7438 ? 7'h7f : 7'h0;
  assign T7438 = T4617[4'h9];
  assign T4618 = T4555 & T4619;
  assign T4619 = 4'h7 == T4554;
  assign T4620 = T4625 | T7439;
  assign T7439 = {T7441, T4621};
  assign T4621 = T7440 & T4622;
  assign T4622 = 9'h80;
  assign T7440 = T4623 ? 9'h1ff : 9'h0;
  assign T4623 = T4624;
  assign T4624 = 1'h1;
  assign T7441 = T7442 ? 8'hff : 8'h0;
  assign T7442 = T4621[4'h8];
  assign T4625 = T4537 & T7443;
  assign T7443 = {T7444, T4626};
  assign T4626 = ~ T4622;
  assign T7444 = T7445 ? 8'hff : 8'h0;
  assign T7445 = T4626[4'h8];
  assign T4627 = T4555 & T4628;
  assign T4628 = 4'h8 == T4554;
  assign T4629 = T4634 | T7446;
  assign T7446 = {T7448, T4630};
  assign T4630 = T7447 & T4631;
  assign T4631 = 8'h40;
  assign T7447 = T4632 ? 8'hff : 8'h0;
  assign T4632 = T4633;
  assign T4633 = 1'h1;
  assign T7448 = T7449 ? 9'h1ff : 9'h0;
  assign T7449 = T4630[3'h7];
  assign T4634 = T4536 & T7450;
  assign T7450 = {T7451, T4635};
  assign T4635 = ~ T4631;
  assign T7451 = T7452 ? 9'h1ff : 9'h0;
  assign T7452 = T4635[3'h7];
  assign T4636 = T4555 & T4637;
  assign T4637 = 4'h9 == T4554;
  assign T4638 = T4643 | T7453;
  assign T7453 = {T7455, T4639};
  assign T4639 = T7454 & T4640;
  assign T4640 = 7'h20;
  assign T7454 = T4641 ? 7'h7f : 7'h0;
  assign T4641 = T4642;
  assign T4642 = 1'h1;
  assign T7455 = T7456 ? 10'h3ff : 10'h0;
  assign T7456 = T4639[3'h6];
  assign T4643 = T4535 & T7457;
  assign T7457 = {T7458, T4644};
  assign T4644 = ~ T4640;
  assign T7458 = T7459 ? 10'h3ff : 10'h0;
  assign T7459 = T4644[3'h6];
  assign T4645 = T4555 & T4646;
  assign T4646 = 4'ha == T4554;
  assign T4647 = T4652 | T7460;
  assign T7460 = {T7462, T4648};
  assign T4648 = T7461 & T4649;
  assign T4649 = 6'h10;
  assign T7461 = T4650 ? 6'h3f : 6'h0;
  assign T4650 = T4651;
  assign T4651 = 1'h1;
  assign T7462 = T7463 ? 11'h7ff : 11'h0;
  assign T7463 = T4648[3'h5];
  assign T4652 = T4534 & T7464;
  assign T7464 = {T7465, T4653};
  assign T4653 = ~ T4649;
  assign T7465 = T7466 ? 11'h7ff : 11'h0;
  assign T7466 = T4653[3'h5];
  assign T4654 = T4555 & T4655;
  assign T4655 = 4'hb == T4554;
  assign T4656 = T4661 | T7467;
  assign T7467 = {T7469, T4657};
  assign T4657 = T7468 & T4658;
  assign T4658 = 5'h8;
  assign T7468 = T4659 ? 5'h1f : 5'h0;
  assign T4659 = T4660;
  assign T4660 = 1'h1;
  assign T7469 = T7470 ? 12'hfff : 12'h0;
  assign T7470 = T4657[3'h4];
  assign T4661 = T4533 & T7471;
  assign T7471 = {T7472, T4662};
  assign T4662 = ~ T4658;
  assign T7472 = T7473 ? 12'hfff : 12'h0;
  assign T7473 = T4662[3'h4];
  assign T4663 = T4555 & T4664;
  assign T4664 = 4'hc == T4554;
  assign T4665 = T4670 | T7474;
  assign T7474 = {T7476, T4666};
  assign T4666 = T7475 & T4667;
  assign T4667 = 4'h4;
  assign T7475 = T4668 ? 4'hf : 4'h0;
  assign T4668 = T4669;
  assign T4669 = 1'h1;
  assign T7476 = T7477 ? 13'h1fff : 13'h0;
  assign T7477 = T4666[2'h3];
  assign T4670 = T4532 & T7478;
  assign T7478 = {T7479, T4671};
  assign T4671 = ~ T4667;
  assign T7479 = T7480 ? 13'h1fff : 13'h0;
  assign T7480 = T4671[2'h3];
  assign T4672 = T4555 & T4673;
  assign T4673 = 4'hd == T4554;
  assign T4674 = T4679 | T7481;
  assign T7481 = {T7483, T4675};
  assign T4675 = T7482 & T4676;
  assign T4676 = 3'h2;
  assign T7482 = T4677 ? 3'h7 : 3'h0;
  assign T4677 = T4678;
  assign T4678 = 1'h1;
  assign T7483 = T7484 ? 14'h3fff : 14'h0;
  assign T7484 = T4675[2'h2];
  assign T4679 = T4531 & T7485;
  assign T7485 = {T7486, T4680};
  assign T4680 = ~ T4676;
  assign T7486 = T7487 ? 14'h3fff : 14'h0;
  assign T7487 = T4680[2'h2];
  assign T4681 = T4555 & T4682;
  assign T4682 = 4'he == T4554;
  assign T4683 = T4688 | T7488;
  assign T7488 = {T7490, T4684};
  assign T4684 = T7489 & T4685;
  assign T4685 = 2'h1;
  assign T7489 = T4686 ? 2'h3 : 2'h0;
  assign T4686 = T4687;
  assign T4687 = 1'h1;
  assign T7490 = T7491 ? 15'h7fff : 15'h0;
  assign T7491 = T4684[1'h1];
  assign T4688 = T4530 & T7492;
  assign T7492 = {T7493, T4689};
  assign T4689 = ~ T4685;
  assign T7493 = T7494 ? 15'h7fff : 15'h0;
  assign T7494 = T4689[1'h1];
  assign T4690 = T4555 & T4691;
  assign T4691 = 4'hf == T4554;
  assign io_V_wire_en_21 = V_wire_en_21;
  assign V_wire_en_21 = T7495;
  assign T7495 = T4692[4'hf:1'h0];
  assign T4692 = T4853 ? T4846 : T4693;
  assign T4693 = T4844 ? T4837 : T4694;
  assign T4694 = T4835 ? T4828 : T4695;
  assign T4695 = T4826 ? T4819 : T4696;
  assign T4696 = T4817 ? T4810 : T4697;
  assign T4697 = T4808 ? T4801 : T4698;
  assign T4698 = T4799 ? T4792 : T4699;
  assign T4699 = T4790 ? T4783 : T4700;
  assign T4700 = T4781 ? T4774 : T4701;
  assign T4701 = T4772 ? T4765 : T4702;
  assign T4702 = T4763 ? T4756 : T4703;
  assign T4703 = T4754 ? T4747 : T4704;
  assign T4704 = T4745 ? T4738 : T4705;
  assign T4705 = T4736 ? T4729 : T4706;
  assign T4706 = T4727 ? T4720 : T4707;
  assign T4707 = T4715 ? T4708 : 17'h0;
  assign T4708 = T4713 | T4709;
  assign T4709 = T7496 & T4710;
  assign T4710 = 17'h8000;
  assign T7496 = T4711 ? 17'h1ffff : 17'h0;
  assign T4711 = T4712;
  assign T4712 = 1'h1;
  assign T4713 = 17'h0 & T4714;
  assign T4714 = ~ T4710;
  assign T4715 = T4718 & T4716;
  assign T4716 = 4'h0 == T4717;
  assign T4717 = LogicBlockModule_21_io_config_V_out[2'h3:1'h0];
  assign T4718 = T4719;
  assign T4719 = LogicBlockModule_21_io_config_V_out[3'h4];
  assign T4720 = T4725 | T7497;
  assign T7497 = {T7499, T4721};
  assign T4721 = T7498 & T4722;
  assign T4722 = 16'h4000;
  assign T7498 = T4723 ? 16'hffff : 16'h0;
  assign T4723 = T4724;
  assign T4724 = 1'h1;
  assign T7499 = T4721[4'hf];
  assign T4725 = T4707 & T7500;
  assign T7500 = {T7501, T4726};
  assign T4726 = ~ T4722;
  assign T7501 = T4726[4'hf];
  assign T4727 = T4718 & T4728;
  assign T4728 = 4'h1 == T4717;
  assign T4729 = T4734 | T7502;
  assign T7502 = {T7504, T4730};
  assign T4730 = T7503 & T4731;
  assign T4731 = 15'h2000;
  assign T7503 = T4732 ? 15'h7fff : 15'h0;
  assign T4732 = T4733;
  assign T4733 = 1'h1;
  assign T7504 = T7505 ? 2'h3 : 2'h0;
  assign T7505 = T4730[4'he];
  assign T4734 = T4706 & T7506;
  assign T7506 = {T7507, T4735};
  assign T4735 = ~ T4731;
  assign T7507 = T7508 ? 2'h3 : 2'h0;
  assign T7508 = T4735[4'he];
  assign T4736 = T4718 & T4737;
  assign T4737 = 4'h2 == T4717;
  assign T4738 = T4743 | T7509;
  assign T7509 = {T7511, T4739};
  assign T4739 = T7510 & T4740;
  assign T4740 = 14'h1000;
  assign T7510 = T4741 ? 14'h3fff : 14'h0;
  assign T4741 = T4742;
  assign T4742 = 1'h1;
  assign T7511 = T7512 ? 3'h7 : 3'h0;
  assign T7512 = T4739[4'hd];
  assign T4743 = T4705 & T7513;
  assign T7513 = {T7514, T4744};
  assign T4744 = ~ T4740;
  assign T7514 = T7515 ? 3'h7 : 3'h0;
  assign T7515 = T4744[4'hd];
  assign T4745 = T4718 & T4746;
  assign T4746 = 4'h3 == T4717;
  assign T4747 = T4752 | T7516;
  assign T7516 = {T7518, T4748};
  assign T4748 = T7517 & T4749;
  assign T4749 = 13'h800;
  assign T7517 = T4750 ? 13'h1fff : 13'h0;
  assign T4750 = T4751;
  assign T4751 = 1'h1;
  assign T7518 = T7519 ? 4'hf : 4'h0;
  assign T7519 = T4748[4'hc];
  assign T4752 = T4704 & T7520;
  assign T7520 = {T7521, T4753};
  assign T4753 = ~ T4749;
  assign T7521 = T7522 ? 4'hf : 4'h0;
  assign T7522 = T4753[4'hc];
  assign T4754 = T4718 & T4755;
  assign T4755 = 4'h4 == T4717;
  assign T4756 = T4761 | T7523;
  assign T7523 = {T7525, T4757};
  assign T4757 = T7524 & T4758;
  assign T4758 = 12'h400;
  assign T7524 = T4759 ? 12'hfff : 12'h0;
  assign T4759 = T4760;
  assign T4760 = 1'h1;
  assign T7525 = T7526 ? 5'h1f : 5'h0;
  assign T7526 = T4757[4'hb];
  assign T4761 = T4703 & T7527;
  assign T7527 = {T7528, T4762};
  assign T4762 = ~ T4758;
  assign T7528 = T7529 ? 5'h1f : 5'h0;
  assign T7529 = T4762[4'hb];
  assign T4763 = T4718 & T4764;
  assign T4764 = 4'h5 == T4717;
  assign T4765 = T4770 | T7530;
  assign T7530 = {T7532, T4766};
  assign T4766 = T7531 & T4767;
  assign T4767 = 11'h200;
  assign T7531 = T4768 ? 11'h7ff : 11'h0;
  assign T4768 = T4769;
  assign T4769 = 1'h1;
  assign T7532 = T7533 ? 6'h3f : 6'h0;
  assign T7533 = T4766[4'ha];
  assign T4770 = T4702 & T7534;
  assign T7534 = {T7535, T4771};
  assign T4771 = ~ T4767;
  assign T7535 = T7536 ? 6'h3f : 6'h0;
  assign T7536 = T4771[4'ha];
  assign T4772 = T4718 & T4773;
  assign T4773 = 4'h6 == T4717;
  assign T4774 = T4779 | T7537;
  assign T7537 = {T7539, T4775};
  assign T4775 = T7538 & T4776;
  assign T4776 = 10'h100;
  assign T7538 = T4777 ? 10'h3ff : 10'h0;
  assign T4777 = T4778;
  assign T4778 = 1'h1;
  assign T7539 = T7540 ? 7'h7f : 7'h0;
  assign T7540 = T4775[4'h9];
  assign T4779 = T4701 & T7541;
  assign T7541 = {T7542, T4780};
  assign T4780 = ~ T4776;
  assign T7542 = T7543 ? 7'h7f : 7'h0;
  assign T7543 = T4780[4'h9];
  assign T4781 = T4718 & T4782;
  assign T4782 = 4'h7 == T4717;
  assign T4783 = T4788 | T7544;
  assign T7544 = {T7546, T4784};
  assign T4784 = T7545 & T4785;
  assign T4785 = 9'h80;
  assign T7545 = T4786 ? 9'h1ff : 9'h0;
  assign T4786 = T4787;
  assign T4787 = 1'h1;
  assign T7546 = T7547 ? 8'hff : 8'h0;
  assign T7547 = T4784[4'h8];
  assign T4788 = T4700 & T7548;
  assign T7548 = {T7549, T4789};
  assign T4789 = ~ T4785;
  assign T7549 = T7550 ? 8'hff : 8'h0;
  assign T7550 = T4789[4'h8];
  assign T4790 = T4718 & T4791;
  assign T4791 = 4'h8 == T4717;
  assign T4792 = T4797 | T7551;
  assign T7551 = {T7553, T4793};
  assign T4793 = T7552 & T4794;
  assign T4794 = 8'h40;
  assign T7552 = T4795 ? 8'hff : 8'h0;
  assign T4795 = T4796;
  assign T4796 = 1'h1;
  assign T7553 = T7554 ? 9'h1ff : 9'h0;
  assign T7554 = T4793[3'h7];
  assign T4797 = T4699 & T7555;
  assign T7555 = {T7556, T4798};
  assign T4798 = ~ T4794;
  assign T7556 = T7557 ? 9'h1ff : 9'h0;
  assign T7557 = T4798[3'h7];
  assign T4799 = T4718 & T4800;
  assign T4800 = 4'h9 == T4717;
  assign T4801 = T4806 | T7558;
  assign T7558 = {T7560, T4802};
  assign T4802 = T7559 & T4803;
  assign T4803 = 7'h20;
  assign T7559 = T4804 ? 7'h7f : 7'h0;
  assign T4804 = T4805;
  assign T4805 = 1'h1;
  assign T7560 = T7561 ? 10'h3ff : 10'h0;
  assign T7561 = T4802[3'h6];
  assign T4806 = T4698 & T7562;
  assign T7562 = {T7563, T4807};
  assign T4807 = ~ T4803;
  assign T7563 = T7564 ? 10'h3ff : 10'h0;
  assign T7564 = T4807[3'h6];
  assign T4808 = T4718 & T4809;
  assign T4809 = 4'ha == T4717;
  assign T4810 = T4815 | T7565;
  assign T7565 = {T7567, T4811};
  assign T4811 = T7566 & T4812;
  assign T4812 = 6'h10;
  assign T7566 = T4813 ? 6'h3f : 6'h0;
  assign T4813 = T4814;
  assign T4814 = 1'h1;
  assign T7567 = T7568 ? 11'h7ff : 11'h0;
  assign T7568 = T4811[3'h5];
  assign T4815 = T4697 & T7569;
  assign T7569 = {T7570, T4816};
  assign T4816 = ~ T4812;
  assign T7570 = T7571 ? 11'h7ff : 11'h0;
  assign T7571 = T4816[3'h5];
  assign T4817 = T4718 & T4818;
  assign T4818 = 4'hb == T4717;
  assign T4819 = T4824 | T7572;
  assign T7572 = {T7574, T4820};
  assign T4820 = T7573 & T4821;
  assign T4821 = 5'h8;
  assign T7573 = T4822 ? 5'h1f : 5'h0;
  assign T4822 = T4823;
  assign T4823 = 1'h1;
  assign T7574 = T7575 ? 12'hfff : 12'h0;
  assign T7575 = T4820[3'h4];
  assign T4824 = T4696 & T7576;
  assign T7576 = {T7577, T4825};
  assign T4825 = ~ T4821;
  assign T7577 = T7578 ? 12'hfff : 12'h0;
  assign T7578 = T4825[3'h4];
  assign T4826 = T4718 & T4827;
  assign T4827 = 4'hc == T4717;
  assign T4828 = T4833 | T7579;
  assign T7579 = {T7581, T4829};
  assign T4829 = T7580 & T4830;
  assign T4830 = 4'h4;
  assign T7580 = T4831 ? 4'hf : 4'h0;
  assign T4831 = T4832;
  assign T4832 = 1'h1;
  assign T7581 = T7582 ? 13'h1fff : 13'h0;
  assign T7582 = T4829[2'h3];
  assign T4833 = T4695 & T7583;
  assign T7583 = {T7584, T4834};
  assign T4834 = ~ T4830;
  assign T7584 = T7585 ? 13'h1fff : 13'h0;
  assign T7585 = T4834[2'h3];
  assign T4835 = T4718 & T4836;
  assign T4836 = 4'hd == T4717;
  assign T4837 = T4842 | T7586;
  assign T7586 = {T7588, T4838};
  assign T4838 = T7587 & T4839;
  assign T4839 = 3'h2;
  assign T7587 = T4840 ? 3'h7 : 3'h0;
  assign T4840 = T4841;
  assign T4841 = 1'h1;
  assign T7588 = T7589 ? 14'h3fff : 14'h0;
  assign T7589 = T4838[2'h2];
  assign T4842 = T4694 & T7590;
  assign T7590 = {T7591, T4843};
  assign T4843 = ~ T4839;
  assign T7591 = T7592 ? 14'h3fff : 14'h0;
  assign T7592 = T4843[2'h2];
  assign T4844 = T4718 & T4845;
  assign T4845 = 4'he == T4717;
  assign T4846 = T4851 | T7593;
  assign T7593 = {T7595, T4847};
  assign T4847 = T7594 & T4848;
  assign T4848 = 2'h1;
  assign T7594 = T4849 ? 2'h3 : 2'h0;
  assign T4849 = T4850;
  assign T4850 = 1'h1;
  assign T7595 = T7596 ? 15'h7fff : 15'h0;
  assign T7596 = T4847[1'h1];
  assign T4851 = T4693 & T7597;
  assign T7597 = {T7598, T4852};
  assign T4852 = ~ T4848;
  assign T7598 = T7599 ? 15'h7fff : 15'h0;
  assign T7599 = T4852[1'h1];
  assign T4853 = T4718 & T4854;
  assign T4854 = 4'hf == T4717;
  assign io_V_wire_en_22 = V_wire_en_22;
  assign V_wire_en_22 = T7600;
  assign T7600 = T4855[4'hf:1'h0];
  assign T4855 = T5016 ? T5009 : T4856;
  assign T4856 = T5007 ? T5000 : T4857;
  assign T4857 = T4998 ? T4991 : T4858;
  assign T4858 = T4989 ? T4982 : T4859;
  assign T4859 = T4980 ? T4973 : T4860;
  assign T4860 = T4971 ? T4964 : T4861;
  assign T4861 = T4962 ? T4955 : T4862;
  assign T4862 = T4953 ? T4946 : T4863;
  assign T4863 = T4944 ? T4937 : T4864;
  assign T4864 = T4935 ? T4928 : T4865;
  assign T4865 = T4926 ? T4919 : T4866;
  assign T4866 = T4917 ? T4910 : T4867;
  assign T4867 = T4908 ? T4901 : T4868;
  assign T4868 = T4899 ? T4892 : T4869;
  assign T4869 = T4890 ? T4883 : T4870;
  assign T4870 = T4878 ? T4871 : 17'h0;
  assign T4871 = T4876 | T4872;
  assign T4872 = T7601 & T4873;
  assign T4873 = 17'h8000;
  assign T7601 = T4874 ? 17'h1ffff : 17'h0;
  assign T4874 = T4875;
  assign T4875 = 1'h1;
  assign T4876 = 17'h0 & T4877;
  assign T4877 = ~ T4873;
  assign T4878 = T4881 & T4879;
  assign T4879 = 4'h0 == T4880;
  assign T4880 = LogicBlockModule_22_io_config_V_out[2'h3:1'h0];
  assign T4881 = T4882;
  assign T4882 = LogicBlockModule_22_io_config_V_out[3'h4];
  assign T4883 = T4888 | T7602;
  assign T7602 = {T7604, T4884};
  assign T4884 = T7603 & T4885;
  assign T4885 = 16'h4000;
  assign T7603 = T4886 ? 16'hffff : 16'h0;
  assign T4886 = T4887;
  assign T4887 = 1'h1;
  assign T7604 = T4884[4'hf];
  assign T4888 = T4870 & T7605;
  assign T7605 = {T7606, T4889};
  assign T4889 = ~ T4885;
  assign T7606 = T4889[4'hf];
  assign T4890 = T4881 & T4891;
  assign T4891 = 4'h1 == T4880;
  assign T4892 = T4897 | T7607;
  assign T7607 = {T7609, T4893};
  assign T4893 = T7608 & T4894;
  assign T4894 = 15'h2000;
  assign T7608 = T4895 ? 15'h7fff : 15'h0;
  assign T4895 = T4896;
  assign T4896 = 1'h1;
  assign T7609 = T7610 ? 2'h3 : 2'h0;
  assign T7610 = T4893[4'he];
  assign T4897 = T4869 & T7611;
  assign T7611 = {T7612, T4898};
  assign T4898 = ~ T4894;
  assign T7612 = T7613 ? 2'h3 : 2'h0;
  assign T7613 = T4898[4'he];
  assign T4899 = T4881 & T4900;
  assign T4900 = 4'h2 == T4880;
  assign T4901 = T4906 | T7614;
  assign T7614 = {T7616, T4902};
  assign T4902 = T7615 & T4903;
  assign T4903 = 14'h1000;
  assign T7615 = T4904 ? 14'h3fff : 14'h0;
  assign T4904 = T4905;
  assign T4905 = 1'h1;
  assign T7616 = T7617 ? 3'h7 : 3'h0;
  assign T7617 = T4902[4'hd];
  assign T4906 = T4868 & T7618;
  assign T7618 = {T7619, T4907};
  assign T4907 = ~ T4903;
  assign T7619 = T7620 ? 3'h7 : 3'h0;
  assign T7620 = T4907[4'hd];
  assign T4908 = T4881 & T4909;
  assign T4909 = 4'h3 == T4880;
  assign T4910 = T4915 | T7621;
  assign T7621 = {T7623, T4911};
  assign T4911 = T7622 & T4912;
  assign T4912 = 13'h800;
  assign T7622 = T4913 ? 13'h1fff : 13'h0;
  assign T4913 = T4914;
  assign T4914 = 1'h1;
  assign T7623 = T7624 ? 4'hf : 4'h0;
  assign T7624 = T4911[4'hc];
  assign T4915 = T4867 & T7625;
  assign T7625 = {T7626, T4916};
  assign T4916 = ~ T4912;
  assign T7626 = T7627 ? 4'hf : 4'h0;
  assign T7627 = T4916[4'hc];
  assign T4917 = T4881 & T4918;
  assign T4918 = 4'h4 == T4880;
  assign T4919 = T4924 | T7628;
  assign T7628 = {T7630, T4920};
  assign T4920 = T7629 & T4921;
  assign T4921 = 12'h400;
  assign T7629 = T4922 ? 12'hfff : 12'h0;
  assign T4922 = T4923;
  assign T4923 = 1'h1;
  assign T7630 = T7631 ? 5'h1f : 5'h0;
  assign T7631 = T4920[4'hb];
  assign T4924 = T4866 & T7632;
  assign T7632 = {T7633, T4925};
  assign T4925 = ~ T4921;
  assign T7633 = T7634 ? 5'h1f : 5'h0;
  assign T7634 = T4925[4'hb];
  assign T4926 = T4881 & T4927;
  assign T4927 = 4'h5 == T4880;
  assign T4928 = T4933 | T7635;
  assign T7635 = {T7637, T4929};
  assign T4929 = T7636 & T4930;
  assign T4930 = 11'h200;
  assign T7636 = T4931 ? 11'h7ff : 11'h0;
  assign T4931 = T4932;
  assign T4932 = 1'h1;
  assign T7637 = T7638 ? 6'h3f : 6'h0;
  assign T7638 = T4929[4'ha];
  assign T4933 = T4865 & T7639;
  assign T7639 = {T7640, T4934};
  assign T4934 = ~ T4930;
  assign T7640 = T7641 ? 6'h3f : 6'h0;
  assign T7641 = T4934[4'ha];
  assign T4935 = T4881 & T4936;
  assign T4936 = 4'h6 == T4880;
  assign T4937 = T4942 | T7642;
  assign T7642 = {T7644, T4938};
  assign T4938 = T7643 & T4939;
  assign T4939 = 10'h100;
  assign T7643 = T4940 ? 10'h3ff : 10'h0;
  assign T4940 = T4941;
  assign T4941 = 1'h1;
  assign T7644 = T7645 ? 7'h7f : 7'h0;
  assign T7645 = T4938[4'h9];
  assign T4942 = T4864 & T7646;
  assign T7646 = {T7647, T4943};
  assign T4943 = ~ T4939;
  assign T7647 = T7648 ? 7'h7f : 7'h0;
  assign T7648 = T4943[4'h9];
  assign T4944 = T4881 & T4945;
  assign T4945 = 4'h7 == T4880;
  assign T4946 = T4951 | T7649;
  assign T7649 = {T7651, T4947};
  assign T4947 = T7650 & T4948;
  assign T4948 = 9'h80;
  assign T7650 = T4949 ? 9'h1ff : 9'h0;
  assign T4949 = T4950;
  assign T4950 = 1'h1;
  assign T7651 = T7652 ? 8'hff : 8'h0;
  assign T7652 = T4947[4'h8];
  assign T4951 = T4863 & T7653;
  assign T7653 = {T7654, T4952};
  assign T4952 = ~ T4948;
  assign T7654 = T7655 ? 8'hff : 8'h0;
  assign T7655 = T4952[4'h8];
  assign T4953 = T4881 & T4954;
  assign T4954 = 4'h8 == T4880;
  assign T4955 = T4960 | T7656;
  assign T7656 = {T7658, T4956};
  assign T4956 = T7657 & T4957;
  assign T4957 = 8'h40;
  assign T7657 = T4958 ? 8'hff : 8'h0;
  assign T4958 = T4959;
  assign T4959 = 1'h1;
  assign T7658 = T7659 ? 9'h1ff : 9'h0;
  assign T7659 = T4956[3'h7];
  assign T4960 = T4862 & T7660;
  assign T7660 = {T7661, T4961};
  assign T4961 = ~ T4957;
  assign T7661 = T7662 ? 9'h1ff : 9'h0;
  assign T7662 = T4961[3'h7];
  assign T4962 = T4881 & T4963;
  assign T4963 = 4'h9 == T4880;
  assign T4964 = T4969 | T7663;
  assign T7663 = {T7665, T4965};
  assign T4965 = T7664 & T4966;
  assign T4966 = 7'h20;
  assign T7664 = T4967 ? 7'h7f : 7'h0;
  assign T4967 = T4968;
  assign T4968 = 1'h1;
  assign T7665 = T7666 ? 10'h3ff : 10'h0;
  assign T7666 = T4965[3'h6];
  assign T4969 = T4861 & T7667;
  assign T7667 = {T7668, T4970};
  assign T4970 = ~ T4966;
  assign T7668 = T7669 ? 10'h3ff : 10'h0;
  assign T7669 = T4970[3'h6];
  assign T4971 = T4881 & T4972;
  assign T4972 = 4'ha == T4880;
  assign T4973 = T4978 | T7670;
  assign T7670 = {T7672, T4974};
  assign T4974 = T7671 & T4975;
  assign T4975 = 6'h10;
  assign T7671 = T4976 ? 6'h3f : 6'h0;
  assign T4976 = T4977;
  assign T4977 = 1'h1;
  assign T7672 = T7673 ? 11'h7ff : 11'h0;
  assign T7673 = T4974[3'h5];
  assign T4978 = T4860 & T7674;
  assign T7674 = {T7675, T4979};
  assign T4979 = ~ T4975;
  assign T7675 = T7676 ? 11'h7ff : 11'h0;
  assign T7676 = T4979[3'h5];
  assign T4980 = T4881 & T4981;
  assign T4981 = 4'hb == T4880;
  assign T4982 = T4987 | T7677;
  assign T7677 = {T7679, T4983};
  assign T4983 = T7678 & T4984;
  assign T4984 = 5'h8;
  assign T7678 = T4985 ? 5'h1f : 5'h0;
  assign T4985 = T4986;
  assign T4986 = 1'h1;
  assign T7679 = T7680 ? 12'hfff : 12'h0;
  assign T7680 = T4983[3'h4];
  assign T4987 = T4859 & T7681;
  assign T7681 = {T7682, T4988};
  assign T4988 = ~ T4984;
  assign T7682 = T7683 ? 12'hfff : 12'h0;
  assign T7683 = T4988[3'h4];
  assign T4989 = T4881 & T4990;
  assign T4990 = 4'hc == T4880;
  assign T4991 = T4996 | T7684;
  assign T7684 = {T7686, T4992};
  assign T4992 = T7685 & T4993;
  assign T4993 = 4'h4;
  assign T7685 = T4994 ? 4'hf : 4'h0;
  assign T4994 = T4995;
  assign T4995 = 1'h1;
  assign T7686 = T7687 ? 13'h1fff : 13'h0;
  assign T7687 = T4992[2'h3];
  assign T4996 = T4858 & T7688;
  assign T7688 = {T7689, T4997};
  assign T4997 = ~ T4993;
  assign T7689 = T7690 ? 13'h1fff : 13'h0;
  assign T7690 = T4997[2'h3];
  assign T4998 = T4881 & T4999;
  assign T4999 = 4'hd == T4880;
  assign T5000 = T5005 | T7691;
  assign T7691 = {T7693, T5001};
  assign T5001 = T7692 & T5002;
  assign T5002 = 3'h2;
  assign T7692 = T5003 ? 3'h7 : 3'h0;
  assign T5003 = T5004;
  assign T5004 = 1'h1;
  assign T7693 = T7694 ? 14'h3fff : 14'h0;
  assign T7694 = T5001[2'h2];
  assign T5005 = T4857 & T7695;
  assign T7695 = {T7696, T5006};
  assign T5006 = ~ T5002;
  assign T7696 = T7697 ? 14'h3fff : 14'h0;
  assign T7697 = T5006[2'h2];
  assign T5007 = T4881 & T5008;
  assign T5008 = 4'he == T4880;
  assign T5009 = T5014 | T7698;
  assign T7698 = {T7700, T5010};
  assign T5010 = T7699 & T5011;
  assign T5011 = 2'h1;
  assign T7699 = T5012 ? 2'h3 : 2'h0;
  assign T5012 = T5013;
  assign T5013 = 1'h1;
  assign T7700 = T7701 ? 15'h7fff : 15'h0;
  assign T7701 = T5010[1'h1];
  assign T5014 = T4856 & T7702;
  assign T7702 = {T7703, T5015};
  assign T5015 = ~ T5011;
  assign T7703 = T7704 ? 15'h7fff : 15'h0;
  assign T7704 = T5015[1'h1];
  assign T5016 = T4881 & T5017;
  assign T5017 = 4'hf == T4880;
  assign io_V_wire_out_0 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_1 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_2 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_3 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_4 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_5 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_6 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_7 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_8 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_9 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_10 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_11 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_12 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_13 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_14 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_15 = LogicBlockModule_io_V_wire_out;
  assign io_V_wire_out_16 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_17 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_18 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_19 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_20 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_21 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_22 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_23 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_24 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_25 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_26 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_27 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_28 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_29 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_30 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_31 = LogicBlockModule_1_io_V_wire_out;
  assign io_V_wire_out_32 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_33 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_34 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_35 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_36 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_37 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_38 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_39 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_40 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_41 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_42 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_43 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_44 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_45 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_46 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_47 = LogicBlockModule_2_io_V_wire_out;
  assign io_V_wire_out_48 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_49 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_50 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_51 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_52 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_53 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_54 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_55 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_56 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_57 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_58 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_59 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_60 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_61 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_62 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_63 = LogicBlockModule_3_io_V_wire_out;
  assign io_V_wire_out_64 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_65 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_66 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_67 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_68 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_69 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_70 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_71 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_72 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_73 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_74 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_75 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_76 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_77 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_78 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_79 = LogicBlockModule_4_io_V_wire_out;
  assign io_V_wire_out_80 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_81 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_82 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_83 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_84 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_85 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_86 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_87 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_88 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_89 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_90 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_91 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_92 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_93 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_94 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_95 = LogicBlockModule_5_io_V_wire_out;
  assign io_V_wire_out_96 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_97 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_98 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_99 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_100 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_101 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_102 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_103 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_104 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_105 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_106 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_107 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_108 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_109 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_110 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_111 = LogicBlockModule_6_io_V_wire_out;
  assign io_V_wire_out_112 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_113 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_114 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_115 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_116 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_117 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_118 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_119 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_120 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_121 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_122 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_123 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_124 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_125 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_126 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_127 = LogicBlockModule_7_io_V_wire_out;
  assign io_V_wire_out_128 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_129 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_130 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_131 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_132 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_133 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_134 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_135 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_136 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_137 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_138 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_139 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_140 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_141 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_142 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_143 = LogicBlockModule_8_io_V_wire_out;
  assign io_V_wire_out_144 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_145 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_146 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_147 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_148 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_149 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_150 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_151 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_152 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_153 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_154 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_155 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_156 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_157 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_158 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_159 = LogicBlockModule_9_io_V_wire_out;
  assign io_V_wire_out_160 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_161 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_162 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_163 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_164 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_165 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_166 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_167 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_168 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_169 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_170 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_171 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_172 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_173 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_174 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_175 = LogicBlockModule_10_io_V_wire_out;
  assign io_V_wire_out_176 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_177 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_178 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_179 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_180 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_181 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_182 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_183 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_184 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_185 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_186 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_187 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_188 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_189 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_190 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_191 = LogicBlockModule_11_io_V_wire_out;
  assign io_V_wire_out_192 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_193 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_194 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_195 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_196 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_197 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_198 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_199 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_200 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_201 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_202 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_203 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_204 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_205 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_206 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_207 = LogicBlockModule_12_io_V_wire_out;
  assign io_V_wire_out_208 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_209 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_210 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_211 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_212 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_213 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_214 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_215 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_216 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_217 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_218 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_219 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_220 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_221 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_222 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_223 = LogicBlockModule_13_io_V_wire_out;
  assign io_V_wire_out_224 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_225 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_226 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_227 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_228 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_229 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_230 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_231 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_232 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_233 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_234 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_235 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_236 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_237 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_238 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_239 = LogicBlockModule_14_io_V_wire_out;
  assign io_V_wire_out_240 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_241 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_242 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_243 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_244 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_245 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_246 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_247 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_248 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_249 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_250 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_251 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_252 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_253 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_254 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_255 = LogicBlockModule_15_io_V_wire_out;
  assign io_V_wire_out_256 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_257 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_258 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_259 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_260 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_261 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_262 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_263 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_264 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_265 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_266 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_267 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_268 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_269 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_270 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_271 = LogicBlockModule_16_io_V_wire_out;
  assign io_V_wire_out_272 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_273 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_274 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_275 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_276 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_277 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_278 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_279 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_280 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_281 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_282 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_283 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_284 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_285 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_286 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_287 = LogicBlockModule_17_io_V_wire_out;
  assign io_V_wire_out_288 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_289 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_290 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_291 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_292 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_293 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_294 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_295 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_296 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_297 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_298 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_299 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_300 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_301 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_302 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_303 = LogicBlockModule_18_io_V_wire_out;
  assign io_V_wire_out_304 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_305 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_306 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_307 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_308 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_309 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_310 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_311 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_312 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_313 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_314 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_315 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_316 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_317 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_318 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_319 = LogicBlockModule_19_io_V_wire_out;
  assign io_V_wire_out_320 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_321 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_322 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_323 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_324 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_325 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_326 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_327 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_328 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_329 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_330 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_331 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_332 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_333 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_334 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_335 = LogicBlockModule_20_io_V_wire_out;
  assign io_V_wire_out_336 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_337 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_338 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_339 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_340 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_341 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_342 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_343 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_344 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_345 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_346 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_347 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_348 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_349 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_350 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_351 = LogicBlockModule_21_io_V_wire_out;
  assign io_V_wire_out_352 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_353 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_354 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_355 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_356 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_357 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_358 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_359 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_360 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_361 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_362 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_363 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_364 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_365 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_366 = LogicBlockModule_22_io_V_wire_out;
  assign io_V_wire_out_367 = LogicBlockModule_22_io_V_wire_out;
  ConfigurationModule ConfigurationModule(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_0 ),
       .io_en( T1268 ),
       .io_out( ConfigurationModule_io_out )
  );
  ConfigurationModule ConfigurationModule_1(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_1 ),
       .io_en( T1267 ),
       .io_out( ConfigurationModule_1_io_out )
  );
  ConfigurationModule ConfigurationModule_2(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_2 ),
       .io_en( T1266 ),
       .io_out( ConfigurationModule_2_io_out )
  );
  ConfigurationModule ConfigurationModule_3(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_3 ),
       .io_en( T1265 ),
       .io_out( ConfigurationModule_3_io_out )
  );
  ConfigurationModule ConfigurationModule_4(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_4 ),
       .io_en( T1264 ),
       .io_out( ConfigurationModule_4_io_out )
  );
  ConfigurationModule ConfigurationModule_5(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_5 ),
       .io_en( T1263 ),
       .io_out( ConfigurationModule_5_io_out )
  );
  ConfigurationModule ConfigurationModule_6(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_6 ),
       .io_en( T1262 ),
       .io_out( ConfigurationModule_6_io_out )
  );
  ConfigurationModule ConfigurationModule_7(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_7 ),
       .io_en( T1261 ),
       .io_out( ConfigurationModule_7_io_out )
  );
  ConfigurationModule ConfigurationModule_8(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_8 ),
       .io_en( T1260 ),
       .io_out( ConfigurationModule_8_io_out )
  );
  ConfigurationModule ConfigurationModule_9(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_9 ),
       .io_en( T1259 ),
       .io_out( ConfigurationModule_9_io_out )
  );
  ConfigurationModule ConfigurationModule_10(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_10 ),
       .io_en( T1258 ),
       .io_out( ConfigurationModule_10_io_out )
  );
  ConfigurationModule ConfigurationModule_11(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_11 ),
       .io_en( T1257 ),
       .io_out( ConfigurationModule_11_io_out )
  );
  ConfigurationModule ConfigurationModule_12(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_12 ),
       .io_en( T1256 ),
       .io_out( ConfigurationModule_12_io_out )
  );
  ConfigurationModule ConfigurationModule_13(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_13 ),
       .io_en( T1255 ),
       .io_out( ConfigurationModule_13_io_out )
  );
  ConfigurationModule ConfigurationModule_14(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_14 ),
       .io_en( T1254 ),
       .io_out( ConfigurationModule_14_io_out )
  );
  ConfigurationModule ConfigurationModule_15(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_15 ),
       .io_en( T1253 ),
       .io_out( ConfigurationModule_15_io_out )
  );
  ConfigurationModule ConfigurationModule_16(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_16 ),
       .io_en( T1252 ),
       .io_out( ConfigurationModule_16_io_out )
  );
  ConfigurationModule ConfigurationModule_17(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_17 ),
       .io_en( T1251 ),
       .io_out( ConfigurationModule_17_io_out )
  );
  ConfigurationModule ConfigurationModule_18(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_18 ),
       .io_en( T1250 ),
       .io_out( ConfigurationModule_18_io_out )
  );
  ConfigurationModule ConfigurationModule_19(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_19 ),
       .io_en( T1249 ),
       .io_out( ConfigurationModule_19_io_out )
  );
  ConfigurationModule ConfigurationModule_20(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_20 ),
       .io_en( T1248 ),
       .io_out( ConfigurationModule_20_io_out )
  );
  ConfigurationModule ConfigurationModule_21(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_21 ),
       .io_en( T1247 ),
       .io_out( ConfigurationModule_21_io_out )
  );
  ConfigurationModule ConfigurationModule_22(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_22 ),
       .io_en( T1246 ),
       .io_out( ConfigurationModule_22_io_out )
  );
  ConfigurationModule ConfigurationModule_23(.clk(clk), .reset(reset),
       .io_in( io_mem_bus_in_23 ),
       .io_en( T1245 ),
       .io_out( ConfigurationModule_23_io_out )
  );
  ControlBlockModule ControlBlockModule(.clk(clk), .reset(reset),
       .io_H_wire_above_in_8( io_H_wire_above_9 ),
       .io_H_wire_above_in_7( io_H_wire_above_8 ),
       .io_H_wire_above_in_6( io_H_wire_above_7 ),
       .io_H_wire_above_in_5( io_H_wire_above_6 ),
       .io_H_wire_above_in_4( io_H_wire_above_5 ),
       .io_H_wire_above_in_3( io_H_wire_above_4 ),
       .io_H_wire_above_in_2( io_H_wire_above_3 ),
       .io_H_wire_above_in_1( io_H_wire_above_2 ),
       .io_H_wire_above_in_0( io_H_wire_above_1 ),
       .io_H_wire_below_in_8( H_wire_below_9 ),
       .io_H_wire_below_in_7( H_wire_below_8 ),
       .io_H_wire_below_in_6( H_wire_below_7 ),
       .io_H_wire_below_in_5( H_wire_below_6 ),
       .io_H_wire_below_in_4( H_wire_below_5 ),
       .io_H_wire_below_in_3( H_wire_below_4 ),
       .io_H_wire_below_in_2( H_wire_below_3 ),
       .io_H_wire_below_in_1( H_wire_below_2 ),
       .io_H_wire_below_in_0( H_wire_below_1 ),
       .io_config( config_23 ),
       .io_Hdir( ControlBlockModule_io_Hdir ),
       //.io_read_demand_access(  )
       //.io_write_demand_access(  )
       //.io_prefetch_demand_access(  )
       //.io_load_transfer_access(  )
       .io_store_transfer_access( ControlBlockModule_io_store_transfer_access ),
       .io_mem_D_or_Z( ControlBlockModule_io_mem_D_or_Z )
  );
  LogicBlockModule LogicBlockModule(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_15 ),
       .io_V_wire_in_14( io_V_wire_in_14 ),
       .io_V_wire_in_13( io_V_wire_in_13 ),
       .io_V_wire_in_12( io_V_wire_in_12 ),
       .io_V_wire_in_11( io_V_wire_in_11 ),
       .io_V_wire_in_10( io_V_wire_in_10 ),
       .io_V_wire_in_9( io_V_wire_in_9 ),
       .io_V_wire_in_8( io_V_wire_in_8 ),
       .io_V_wire_in_7( io_V_wire_in_7 ),
       .io_V_wire_in_6( io_V_wire_in_6 ),
       .io_V_wire_in_5( io_V_wire_in_5 ),
       .io_V_wire_in_4( io_V_wire_in_4 ),
       .io_V_wire_in_3( io_V_wire_in_3 ),
       .io_V_wire_in_2( io_V_wire_in_2 ),
       .io_V_wire_in_1( io_V_wire_in_1 ),
       .io_V_wire_in_0( io_V_wire_in_0 ),
       .io_H_wire_above_in_10( io_H_wire_above_32 ),
       .io_H_wire_above_in_9( io_H_wire_above_31 ),
       .io_H_wire_above_in_8( io_H_wire_above_30 ),
       .io_H_wire_above_in_7( io_H_wire_above_29 ),
       .io_H_wire_above_in_6( io_H_wire_above_28 ),
       .io_H_wire_above_in_5( io_H_wire_above_27 ),
       .io_H_wire_above_in_4( io_H_wire_above_26 ),
       .io_H_wire_above_in_3( io_H_wire_above_25 ),
       .io_H_wire_above_in_2( io_H_wire_above_24 ),
       .io_H_wire_above_in_1( io_H_wire_above_23 ),
       .io_H_wire_above_in_0( io_H_wire_above_22 ),
       .io_H_wire_below_in_10( H_wire_below_32 ),
       .io_H_wire_below_in_9( H_wire_below_31 ),
       .io_H_wire_below_in_8( H_wire_below_30 ),
       .io_H_wire_below_in_7( H_wire_below_29 ),
       .io_H_wire_below_in_6( H_wire_below_28 ),
       .io_H_wire_below_in_5( H_wire_below_27 ),
       .io_H_wire_below_in_4( H_wire_below_26 ),
       .io_H_wire_below_in_3( H_wire_below_25 ),
       .io_H_wire_below_in_2( H_wire_below_24 ),
       .io_H_wire_below_in_1( H_wire_below_23 ),
       .io_H_wire_below_in_0( H_wire_below_22 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_0 ),
       .io_shift_X_in_2( 1'h0 ),
       .io_shift_X_in_1( 1'h0 ),
       .io_shift_X_in_0( 1'h0 ),
       .io_H_out_above( io_H_out_above_0 ),
       .io_shift_carry_in( 1'h0 ),
       .io_carry_in( 1'h0 ),
       .io_shift_X_out_2( LogicBlockModule_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_io_carry_out ),
       .io_store_en( T1242 ),
       .io_mem_D_or_Z( T1237 ),
       .io_config( config_0 ),
       .io_mem_bus_out( LogicBlockModule_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_1(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_31 ),
       .io_V_wire_in_14( io_V_wire_in_30 ),
       .io_V_wire_in_13( io_V_wire_in_29 ),
       .io_V_wire_in_12( io_V_wire_in_28 ),
       .io_V_wire_in_11( io_V_wire_in_27 ),
       .io_V_wire_in_10( io_V_wire_in_26 ),
       .io_V_wire_in_9( io_V_wire_in_25 ),
       .io_V_wire_in_8( io_V_wire_in_24 ),
       .io_V_wire_in_7( io_V_wire_in_23 ),
       .io_V_wire_in_6( io_V_wire_in_22 ),
       .io_V_wire_in_5( io_V_wire_in_21 ),
       .io_V_wire_in_4( io_V_wire_in_20 ),
       .io_V_wire_in_3( io_V_wire_in_19 ),
       .io_V_wire_in_2( io_V_wire_in_18 ),
       .io_V_wire_in_1( io_V_wire_in_17 ),
       .io_V_wire_in_0( io_V_wire_in_16 ),
       .io_H_wire_above_in_10( io_H_wire_above_31 ),
       .io_H_wire_above_in_9( io_H_wire_above_30 ),
       .io_H_wire_above_in_8( io_H_wire_above_29 ),
       .io_H_wire_above_in_7( io_H_wire_above_28 ),
       .io_H_wire_above_in_6( io_H_wire_above_27 ),
       .io_H_wire_above_in_5( io_H_wire_above_26 ),
       .io_H_wire_above_in_4( io_H_wire_above_25 ),
       .io_H_wire_above_in_3( io_H_wire_above_24 ),
       .io_H_wire_above_in_2( io_H_wire_above_23 ),
       .io_H_wire_above_in_1( io_H_wire_above_22 ),
       .io_H_wire_above_in_0( io_H_wire_above_21 ),
       .io_H_wire_below_in_10( H_wire_below_31 ),
       .io_H_wire_below_in_9( H_wire_below_30 ),
       .io_H_wire_below_in_8( H_wire_below_29 ),
       .io_H_wire_below_in_7( H_wire_below_28 ),
       .io_H_wire_below_in_6( H_wire_below_27 ),
       .io_H_wire_below_in_5( H_wire_below_26 ),
       .io_H_wire_below_in_4( H_wire_below_25 ),
       .io_H_wire_below_in_3( H_wire_below_24 ),
       .io_H_wire_below_in_2( H_wire_below_23 ),
       .io_H_wire_below_in_1( H_wire_below_22 ),
       .io_H_wire_below_in_0( H_wire_below_21 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_1 ),
       .io_shift_X_in_2( LogicBlockModule_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_1 ),
       .io_shift_carry_in( LogicBlockModule_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_1_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_1_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_1_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_1_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_1_io_carry_out ),
       .io_store_en( T1234 ),
       .io_mem_D_or_Z( T1229 ),
       .io_config( config_1 ),
       .io_mem_bus_out( LogicBlockModule_1_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_1_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_1_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_1_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_1_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_1_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_2(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_47 ),
       .io_V_wire_in_14( io_V_wire_in_46 ),
       .io_V_wire_in_13( io_V_wire_in_45 ),
       .io_V_wire_in_12( io_V_wire_in_44 ),
       .io_V_wire_in_11( io_V_wire_in_43 ),
       .io_V_wire_in_10( io_V_wire_in_42 ),
       .io_V_wire_in_9( io_V_wire_in_41 ),
       .io_V_wire_in_8( io_V_wire_in_40 ),
       .io_V_wire_in_7( io_V_wire_in_39 ),
       .io_V_wire_in_6( io_V_wire_in_38 ),
       .io_V_wire_in_5( io_V_wire_in_37 ),
       .io_V_wire_in_4( io_V_wire_in_36 ),
       .io_V_wire_in_3( io_V_wire_in_35 ),
       .io_V_wire_in_2( io_V_wire_in_34 ),
       .io_V_wire_in_1( io_V_wire_in_33 ),
       .io_V_wire_in_0( io_V_wire_in_32 ),
       .io_H_wire_above_in_10( io_H_wire_above_30 ),
       .io_H_wire_above_in_9( io_H_wire_above_29 ),
       .io_H_wire_above_in_8( io_H_wire_above_28 ),
       .io_H_wire_above_in_7( io_H_wire_above_27 ),
       .io_H_wire_above_in_6( io_H_wire_above_26 ),
       .io_H_wire_above_in_5( io_H_wire_above_25 ),
       .io_H_wire_above_in_4( io_H_wire_above_24 ),
       .io_H_wire_above_in_3( io_H_wire_above_23 ),
       .io_H_wire_above_in_2( io_H_wire_above_22 ),
       .io_H_wire_above_in_1( io_H_wire_above_21 ),
       .io_H_wire_above_in_0( io_H_wire_above_20 ),
       .io_H_wire_below_in_10( H_wire_below_30 ),
       .io_H_wire_below_in_9( H_wire_below_29 ),
       .io_H_wire_below_in_8( H_wire_below_28 ),
       .io_H_wire_below_in_7( H_wire_below_27 ),
       .io_H_wire_below_in_6( H_wire_below_26 ),
       .io_H_wire_below_in_5( H_wire_below_25 ),
       .io_H_wire_below_in_4( H_wire_below_24 ),
       .io_H_wire_below_in_3( H_wire_below_23 ),
       .io_H_wire_below_in_2( H_wire_below_22 ),
       .io_H_wire_below_in_1( H_wire_below_21 ),
       .io_H_wire_below_in_0( H_wire_below_20 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_2 ),
       .io_shift_X_in_2( LogicBlockModule_1_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_1_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_1_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_2 ),
       .io_shift_carry_in( LogicBlockModule_1_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_1_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_2_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_2_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_2_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_2_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_2_io_carry_out ),
       .io_store_en( T1226 ),
       .io_mem_D_or_Z( T1221 ),
       .io_config( config_2 ),
       .io_mem_bus_out( LogicBlockModule_2_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_2_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_2_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_2_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_2_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_2_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_3(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_63 ),
       .io_V_wire_in_14( io_V_wire_in_62 ),
       .io_V_wire_in_13( io_V_wire_in_61 ),
       .io_V_wire_in_12( io_V_wire_in_60 ),
       .io_V_wire_in_11( io_V_wire_in_59 ),
       .io_V_wire_in_10( io_V_wire_in_58 ),
       .io_V_wire_in_9( io_V_wire_in_57 ),
       .io_V_wire_in_8( io_V_wire_in_56 ),
       .io_V_wire_in_7( io_V_wire_in_55 ),
       .io_V_wire_in_6( io_V_wire_in_54 ),
       .io_V_wire_in_5( io_V_wire_in_53 ),
       .io_V_wire_in_4( io_V_wire_in_52 ),
       .io_V_wire_in_3( io_V_wire_in_51 ),
       .io_V_wire_in_2( io_V_wire_in_50 ),
       .io_V_wire_in_1( io_V_wire_in_49 ),
       .io_V_wire_in_0( io_V_wire_in_48 ),
       .io_H_wire_above_in_10( io_H_wire_above_29 ),
       .io_H_wire_above_in_9( io_H_wire_above_28 ),
       .io_H_wire_above_in_8( io_H_wire_above_27 ),
       .io_H_wire_above_in_7( io_H_wire_above_26 ),
       .io_H_wire_above_in_6( io_H_wire_above_25 ),
       .io_H_wire_above_in_5( io_H_wire_above_24 ),
       .io_H_wire_above_in_4( io_H_wire_above_23 ),
       .io_H_wire_above_in_3( io_H_wire_above_22 ),
       .io_H_wire_above_in_2( io_H_wire_above_21 ),
       .io_H_wire_above_in_1( io_H_wire_above_20 ),
       .io_H_wire_above_in_0( io_H_wire_above_19 ),
       .io_H_wire_below_in_10( H_wire_below_29 ),
       .io_H_wire_below_in_9( H_wire_below_28 ),
       .io_H_wire_below_in_8( H_wire_below_27 ),
       .io_H_wire_below_in_7( H_wire_below_26 ),
       .io_H_wire_below_in_6( H_wire_below_25 ),
       .io_H_wire_below_in_5( H_wire_below_24 ),
       .io_H_wire_below_in_4( H_wire_below_23 ),
       .io_H_wire_below_in_3( H_wire_below_22 ),
       .io_H_wire_below_in_2( H_wire_below_21 ),
       .io_H_wire_below_in_1( H_wire_below_20 ),
       .io_H_wire_below_in_0( H_wire_below_19 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_3 ),
       .io_shift_X_in_2( LogicBlockModule_2_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_2_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_2_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_3 ),
       .io_shift_carry_in( LogicBlockModule_2_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_2_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_3_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_3_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_3_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_3_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_3_io_carry_out ),
       .io_store_en( T1218 ),
       .io_mem_D_or_Z( T1213 ),
       .io_config( config_3 ),
       .io_mem_bus_out( LogicBlockModule_3_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_3_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_3_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_3_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_3_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_3_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_4(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_79 ),
       .io_V_wire_in_14( io_V_wire_in_78 ),
       .io_V_wire_in_13( io_V_wire_in_77 ),
       .io_V_wire_in_12( io_V_wire_in_76 ),
       .io_V_wire_in_11( io_V_wire_in_75 ),
       .io_V_wire_in_10( io_V_wire_in_74 ),
       .io_V_wire_in_9( io_V_wire_in_73 ),
       .io_V_wire_in_8( io_V_wire_in_72 ),
       .io_V_wire_in_7( io_V_wire_in_71 ),
       .io_V_wire_in_6( io_V_wire_in_70 ),
       .io_V_wire_in_5( io_V_wire_in_69 ),
       .io_V_wire_in_4( io_V_wire_in_68 ),
       .io_V_wire_in_3( io_V_wire_in_67 ),
       .io_V_wire_in_2( io_V_wire_in_66 ),
       .io_V_wire_in_1( io_V_wire_in_65 ),
       .io_V_wire_in_0( io_V_wire_in_64 ),
       .io_H_wire_above_in_10( io_H_wire_above_28 ),
       .io_H_wire_above_in_9( io_H_wire_above_27 ),
       .io_H_wire_above_in_8( io_H_wire_above_26 ),
       .io_H_wire_above_in_7( io_H_wire_above_25 ),
       .io_H_wire_above_in_6( io_H_wire_above_24 ),
       .io_H_wire_above_in_5( io_H_wire_above_23 ),
       .io_H_wire_above_in_4( io_H_wire_above_22 ),
       .io_H_wire_above_in_3( io_H_wire_above_21 ),
       .io_H_wire_above_in_2( io_H_wire_above_20 ),
       .io_H_wire_above_in_1( io_H_wire_above_19 ),
       .io_H_wire_above_in_0( io_H_wire_above_18 ),
       .io_H_wire_below_in_10( H_wire_below_28 ),
       .io_H_wire_below_in_9( H_wire_below_27 ),
       .io_H_wire_below_in_8( H_wire_below_26 ),
       .io_H_wire_below_in_7( H_wire_below_25 ),
       .io_H_wire_below_in_6( H_wire_below_24 ),
       .io_H_wire_below_in_5( H_wire_below_23 ),
       .io_H_wire_below_in_4( H_wire_below_22 ),
       .io_H_wire_below_in_3( H_wire_below_21 ),
       .io_H_wire_below_in_2( H_wire_below_20 ),
       .io_H_wire_below_in_1( H_wire_below_19 ),
       .io_H_wire_below_in_0( H_wire_below_18 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_4 ),
       .io_shift_X_in_2( LogicBlockModule_3_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_3_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_3_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_4 ),
       .io_shift_carry_in( LogicBlockModule_3_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_3_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_4_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_4_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_4_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_4_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_4_io_carry_out ),
       .io_store_en( T1210 ),
       .io_mem_D_or_Z( T1205 ),
       .io_config( config_4 ),
       .io_mem_bus_out( LogicBlockModule_4_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_4_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_4_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_4_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_4_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_4_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_5(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_95 ),
       .io_V_wire_in_14( io_V_wire_in_94 ),
       .io_V_wire_in_13( io_V_wire_in_93 ),
       .io_V_wire_in_12( io_V_wire_in_92 ),
       .io_V_wire_in_11( io_V_wire_in_91 ),
       .io_V_wire_in_10( io_V_wire_in_90 ),
       .io_V_wire_in_9( io_V_wire_in_89 ),
       .io_V_wire_in_8( io_V_wire_in_88 ),
       .io_V_wire_in_7( io_V_wire_in_87 ),
       .io_V_wire_in_6( io_V_wire_in_86 ),
       .io_V_wire_in_5( io_V_wire_in_85 ),
       .io_V_wire_in_4( io_V_wire_in_84 ),
       .io_V_wire_in_3( io_V_wire_in_83 ),
       .io_V_wire_in_2( io_V_wire_in_82 ),
       .io_V_wire_in_1( io_V_wire_in_81 ),
       .io_V_wire_in_0( io_V_wire_in_80 ),
       .io_H_wire_above_in_10( io_H_wire_above_27 ),
       .io_H_wire_above_in_9( io_H_wire_above_26 ),
       .io_H_wire_above_in_8( io_H_wire_above_25 ),
       .io_H_wire_above_in_7( io_H_wire_above_24 ),
       .io_H_wire_above_in_6( io_H_wire_above_23 ),
       .io_H_wire_above_in_5( io_H_wire_above_22 ),
       .io_H_wire_above_in_4( io_H_wire_above_21 ),
       .io_H_wire_above_in_3( io_H_wire_above_20 ),
       .io_H_wire_above_in_2( io_H_wire_above_19 ),
       .io_H_wire_above_in_1( io_H_wire_above_18 ),
       .io_H_wire_above_in_0( io_H_wire_above_17 ),
       .io_H_wire_below_in_10( H_wire_below_27 ),
       .io_H_wire_below_in_9( H_wire_below_26 ),
       .io_H_wire_below_in_8( H_wire_below_25 ),
       .io_H_wire_below_in_7( H_wire_below_24 ),
       .io_H_wire_below_in_6( H_wire_below_23 ),
       .io_H_wire_below_in_5( H_wire_below_22 ),
       .io_H_wire_below_in_4( H_wire_below_21 ),
       .io_H_wire_below_in_3( H_wire_below_20 ),
       .io_H_wire_below_in_2( H_wire_below_19 ),
       .io_H_wire_below_in_1( H_wire_below_18 ),
       .io_H_wire_below_in_0( H_wire_below_17 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_5 ),
       .io_shift_X_in_2( LogicBlockModule_4_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_4_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_4_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_5 ),
       .io_shift_carry_in( LogicBlockModule_4_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_4_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_5_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_5_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_5_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_5_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_5_io_carry_out ),
       .io_store_en( T1202 ),
       .io_mem_D_or_Z( T1197 ),
       .io_config( config_5 ),
       .io_mem_bus_out( LogicBlockModule_5_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_5_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_5_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_5_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_5_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_5_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_6(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_111 ),
       .io_V_wire_in_14( io_V_wire_in_110 ),
       .io_V_wire_in_13( io_V_wire_in_109 ),
       .io_V_wire_in_12( io_V_wire_in_108 ),
       .io_V_wire_in_11( io_V_wire_in_107 ),
       .io_V_wire_in_10( io_V_wire_in_106 ),
       .io_V_wire_in_9( io_V_wire_in_105 ),
       .io_V_wire_in_8( io_V_wire_in_104 ),
       .io_V_wire_in_7( io_V_wire_in_103 ),
       .io_V_wire_in_6( io_V_wire_in_102 ),
       .io_V_wire_in_5( io_V_wire_in_101 ),
       .io_V_wire_in_4( io_V_wire_in_100 ),
       .io_V_wire_in_3( io_V_wire_in_99 ),
       .io_V_wire_in_2( io_V_wire_in_98 ),
       .io_V_wire_in_1( io_V_wire_in_97 ),
       .io_V_wire_in_0( io_V_wire_in_96 ),
       .io_H_wire_above_in_10( io_H_wire_above_26 ),
       .io_H_wire_above_in_9( io_H_wire_above_25 ),
       .io_H_wire_above_in_8( io_H_wire_above_24 ),
       .io_H_wire_above_in_7( io_H_wire_above_23 ),
       .io_H_wire_above_in_6( io_H_wire_above_22 ),
       .io_H_wire_above_in_5( io_H_wire_above_21 ),
       .io_H_wire_above_in_4( io_H_wire_above_20 ),
       .io_H_wire_above_in_3( io_H_wire_above_19 ),
       .io_H_wire_above_in_2( io_H_wire_above_18 ),
       .io_H_wire_above_in_1( io_H_wire_above_17 ),
       .io_H_wire_above_in_0( io_H_wire_above_16 ),
       .io_H_wire_below_in_10( H_wire_below_26 ),
       .io_H_wire_below_in_9( H_wire_below_25 ),
       .io_H_wire_below_in_8( H_wire_below_24 ),
       .io_H_wire_below_in_7( H_wire_below_23 ),
       .io_H_wire_below_in_6( H_wire_below_22 ),
       .io_H_wire_below_in_5( H_wire_below_21 ),
       .io_H_wire_below_in_4( H_wire_below_20 ),
       .io_H_wire_below_in_3( H_wire_below_19 ),
       .io_H_wire_below_in_2( H_wire_below_18 ),
       .io_H_wire_below_in_1( H_wire_below_17 ),
       .io_H_wire_below_in_0( H_wire_below_16 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_6 ),
       .io_shift_X_in_2( LogicBlockModule_5_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_5_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_5_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_6 ),
       .io_shift_carry_in( LogicBlockModule_5_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_5_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_6_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_6_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_6_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_6_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_6_io_carry_out ),
       .io_store_en( T1194 ),
       .io_mem_D_or_Z( T1189 ),
       .io_config( config_6 ),
       .io_mem_bus_out( LogicBlockModule_6_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_6_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_6_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_6_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_6_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_6_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_7(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_127 ),
       .io_V_wire_in_14( io_V_wire_in_126 ),
       .io_V_wire_in_13( io_V_wire_in_125 ),
       .io_V_wire_in_12( io_V_wire_in_124 ),
       .io_V_wire_in_11( io_V_wire_in_123 ),
       .io_V_wire_in_10( io_V_wire_in_122 ),
       .io_V_wire_in_9( io_V_wire_in_121 ),
       .io_V_wire_in_8( io_V_wire_in_120 ),
       .io_V_wire_in_7( io_V_wire_in_119 ),
       .io_V_wire_in_6( io_V_wire_in_118 ),
       .io_V_wire_in_5( io_V_wire_in_117 ),
       .io_V_wire_in_4( io_V_wire_in_116 ),
       .io_V_wire_in_3( io_V_wire_in_115 ),
       .io_V_wire_in_2( io_V_wire_in_114 ),
       .io_V_wire_in_1( io_V_wire_in_113 ),
       .io_V_wire_in_0( io_V_wire_in_112 ),
       .io_H_wire_above_in_10( io_H_wire_above_25 ),
       .io_H_wire_above_in_9( io_H_wire_above_24 ),
       .io_H_wire_above_in_8( io_H_wire_above_23 ),
       .io_H_wire_above_in_7( io_H_wire_above_22 ),
       .io_H_wire_above_in_6( io_H_wire_above_21 ),
       .io_H_wire_above_in_5( io_H_wire_above_20 ),
       .io_H_wire_above_in_4( io_H_wire_above_19 ),
       .io_H_wire_above_in_3( io_H_wire_above_18 ),
       .io_H_wire_above_in_2( io_H_wire_above_17 ),
       .io_H_wire_above_in_1( io_H_wire_above_16 ),
       .io_H_wire_above_in_0( io_H_wire_above_15 ),
       .io_H_wire_below_in_10( H_wire_below_25 ),
       .io_H_wire_below_in_9( H_wire_below_24 ),
       .io_H_wire_below_in_8( H_wire_below_23 ),
       .io_H_wire_below_in_7( H_wire_below_22 ),
       .io_H_wire_below_in_6( H_wire_below_21 ),
       .io_H_wire_below_in_5( H_wire_below_20 ),
       .io_H_wire_below_in_4( H_wire_below_19 ),
       .io_H_wire_below_in_3( H_wire_below_18 ),
       .io_H_wire_below_in_2( H_wire_below_17 ),
       .io_H_wire_below_in_1( H_wire_below_16 ),
       .io_H_wire_below_in_0( H_wire_below_15 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_7 ),
       .io_shift_X_in_2( LogicBlockModule_6_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_6_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_6_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_7 ),
       .io_shift_carry_in( LogicBlockModule_6_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_6_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_7_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_7_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_7_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_7_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_7_io_carry_out ),
       .io_store_en( T1186 ),
       .io_mem_D_or_Z( T1181 ),
       .io_config( config_7 ),
       .io_mem_bus_out( LogicBlockModule_7_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_7_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_7_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_7_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_7_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_7_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_8(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_143 ),
       .io_V_wire_in_14( io_V_wire_in_142 ),
       .io_V_wire_in_13( io_V_wire_in_141 ),
       .io_V_wire_in_12( io_V_wire_in_140 ),
       .io_V_wire_in_11( io_V_wire_in_139 ),
       .io_V_wire_in_10( io_V_wire_in_138 ),
       .io_V_wire_in_9( io_V_wire_in_137 ),
       .io_V_wire_in_8( io_V_wire_in_136 ),
       .io_V_wire_in_7( io_V_wire_in_135 ),
       .io_V_wire_in_6( io_V_wire_in_134 ),
       .io_V_wire_in_5( io_V_wire_in_133 ),
       .io_V_wire_in_4( io_V_wire_in_132 ),
       .io_V_wire_in_3( io_V_wire_in_131 ),
       .io_V_wire_in_2( io_V_wire_in_130 ),
       .io_V_wire_in_1( io_V_wire_in_129 ),
       .io_V_wire_in_0( io_V_wire_in_128 ),
       .io_H_wire_above_in_10( io_H_wire_above_24 ),
       .io_H_wire_above_in_9( io_H_wire_above_23 ),
       .io_H_wire_above_in_8( io_H_wire_above_22 ),
       .io_H_wire_above_in_7( io_H_wire_above_21 ),
       .io_H_wire_above_in_6( io_H_wire_above_20 ),
       .io_H_wire_above_in_5( io_H_wire_above_19 ),
       .io_H_wire_above_in_4( io_H_wire_above_18 ),
       .io_H_wire_above_in_3( io_H_wire_above_17 ),
       .io_H_wire_above_in_2( io_H_wire_above_16 ),
       .io_H_wire_above_in_1( io_H_wire_above_15 ),
       .io_H_wire_above_in_0( io_H_wire_above_14 ),
       .io_H_wire_below_in_10( H_wire_below_24 ),
       .io_H_wire_below_in_9( H_wire_below_23 ),
       .io_H_wire_below_in_8( H_wire_below_22 ),
       .io_H_wire_below_in_7( H_wire_below_21 ),
       .io_H_wire_below_in_6( H_wire_below_20 ),
       .io_H_wire_below_in_5( H_wire_below_19 ),
       .io_H_wire_below_in_4( H_wire_below_18 ),
       .io_H_wire_below_in_3( H_wire_below_17 ),
       .io_H_wire_below_in_2( H_wire_below_16 ),
       .io_H_wire_below_in_1( H_wire_below_15 ),
       .io_H_wire_below_in_0( H_wire_below_14 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_8 ),
       .io_shift_X_in_2( LogicBlockModule_7_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_7_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_7_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_8 ),
       .io_shift_carry_in( LogicBlockModule_7_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_7_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_8_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_8_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_8_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_8_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_8_io_carry_out ),
       .io_store_en( T1178 ),
       .io_mem_D_or_Z( T1173 ),
       .io_config( config_8 ),
       .io_mem_bus_out( LogicBlockModule_8_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_8_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_8_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_8_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_8_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_8_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_9(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_159 ),
       .io_V_wire_in_14( io_V_wire_in_158 ),
       .io_V_wire_in_13( io_V_wire_in_157 ),
       .io_V_wire_in_12( io_V_wire_in_156 ),
       .io_V_wire_in_11( io_V_wire_in_155 ),
       .io_V_wire_in_10( io_V_wire_in_154 ),
       .io_V_wire_in_9( io_V_wire_in_153 ),
       .io_V_wire_in_8( io_V_wire_in_152 ),
       .io_V_wire_in_7( io_V_wire_in_151 ),
       .io_V_wire_in_6( io_V_wire_in_150 ),
       .io_V_wire_in_5( io_V_wire_in_149 ),
       .io_V_wire_in_4( io_V_wire_in_148 ),
       .io_V_wire_in_3( io_V_wire_in_147 ),
       .io_V_wire_in_2( io_V_wire_in_146 ),
       .io_V_wire_in_1( io_V_wire_in_145 ),
       .io_V_wire_in_0( io_V_wire_in_144 ),
       .io_H_wire_above_in_10( io_H_wire_above_23 ),
       .io_H_wire_above_in_9( io_H_wire_above_22 ),
       .io_H_wire_above_in_8( io_H_wire_above_21 ),
       .io_H_wire_above_in_7( io_H_wire_above_20 ),
       .io_H_wire_above_in_6( io_H_wire_above_19 ),
       .io_H_wire_above_in_5( io_H_wire_above_18 ),
       .io_H_wire_above_in_4( io_H_wire_above_17 ),
       .io_H_wire_above_in_3( io_H_wire_above_16 ),
       .io_H_wire_above_in_2( io_H_wire_above_15 ),
       .io_H_wire_above_in_1( io_H_wire_above_14 ),
       .io_H_wire_above_in_0( io_H_wire_above_13 ),
       .io_H_wire_below_in_10( H_wire_below_23 ),
       .io_H_wire_below_in_9( H_wire_below_22 ),
       .io_H_wire_below_in_8( H_wire_below_21 ),
       .io_H_wire_below_in_7( H_wire_below_20 ),
       .io_H_wire_below_in_6( H_wire_below_19 ),
       .io_H_wire_below_in_5( H_wire_below_18 ),
       .io_H_wire_below_in_4( H_wire_below_17 ),
       .io_H_wire_below_in_3( H_wire_below_16 ),
       .io_H_wire_below_in_2( H_wire_below_15 ),
       .io_H_wire_below_in_1( H_wire_below_14 ),
       .io_H_wire_below_in_0( H_wire_below_13 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_9 ),
       .io_shift_X_in_2( LogicBlockModule_8_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_8_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_8_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_9 ),
       .io_shift_carry_in( LogicBlockModule_8_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_8_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_9_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_9_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_9_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_9_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_9_io_carry_out ),
       .io_store_en( T1170 ),
       .io_mem_D_or_Z( T1165 ),
       .io_config( config_9 ),
       .io_mem_bus_out( LogicBlockModule_9_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_9_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_9_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_9_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_9_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_9_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_10(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_175 ),
       .io_V_wire_in_14( io_V_wire_in_174 ),
       .io_V_wire_in_13( io_V_wire_in_173 ),
       .io_V_wire_in_12( io_V_wire_in_172 ),
       .io_V_wire_in_11( io_V_wire_in_171 ),
       .io_V_wire_in_10( io_V_wire_in_170 ),
       .io_V_wire_in_9( io_V_wire_in_169 ),
       .io_V_wire_in_8( io_V_wire_in_168 ),
       .io_V_wire_in_7( io_V_wire_in_167 ),
       .io_V_wire_in_6( io_V_wire_in_166 ),
       .io_V_wire_in_5( io_V_wire_in_165 ),
       .io_V_wire_in_4( io_V_wire_in_164 ),
       .io_V_wire_in_3( io_V_wire_in_163 ),
       .io_V_wire_in_2( io_V_wire_in_162 ),
       .io_V_wire_in_1( io_V_wire_in_161 ),
       .io_V_wire_in_0( io_V_wire_in_160 ),
       .io_H_wire_above_in_10( io_H_wire_above_22 ),
       .io_H_wire_above_in_9( io_H_wire_above_21 ),
       .io_H_wire_above_in_8( io_H_wire_above_20 ),
       .io_H_wire_above_in_7( io_H_wire_above_19 ),
       .io_H_wire_above_in_6( io_H_wire_above_18 ),
       .io_H_wire_above_in_5( io_H_wire_above_17 ),
       .io_H_wire_above_in_4( io_H_wire_above_16 ),
       .io_H_wire_above_in_3( io_H_wire_above_15 ),
       .io_H_wire_above_in_2( io_H_wire_above_14 ),
       .io_H_wire_above_in_1( io_H_wire_above_13 ),
       .io_H_wire_above_in_0( io_H_wire_above_12 ),
       .io_H_wire_below_in_10( H_wire_below_22 ),
       .io_H_wire_below_in_9( H_wire_below_21 ),
       .io_H_wire_below_in_8( H_wire_below_20 ),
       .io_H_wire_below_in_7( H_wire_below_19 ),
       .io_H_wire_below_in_6( H_wire_below_18 ),
       .io_H_wire_below_in_5( H_wire_below_17 ),
       .io_H_wire_below_in_4( H_wire_below_16 ),
       .io_H_wire_below_in_3( H_wire_below_15 ),
       .io_H_wire_below_in_2( H_wire_below_14 ),
       .io_H_wire_below_in_1( H_wire_below_13 ),
       .io_H_wire_below_in_0( H_wire_below_12 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_10 ),
       .io_shift_X_in_2( LogicBlockModule_9_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_9_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_9_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_10 ),
       .io_shift_carry_in( LogicBlockModule_9_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_9_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_10_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_10_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_10_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_10_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_10_io_carry_out ),
       .io_store_en( T1162 ),
       .io_mem_D_or_Z( T1157 ),
       .io_config( config_10 ),
       .io_mem_bus_out( LogicBlockModule_10_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_10_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_10_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_10_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_10_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_10_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_11(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_191 ),
       .io_V_wire_in_14( io_V_wire_in_190 ),
       .io_V_wire_in_13( io_V_wire_in_189 ),
       .io_V_wire_in_12( io_V_wire_in_188 ),
       .io_V_wire_in_11( io_V_wire_in_187 ),
       .io_V_wire_in_10( io_V_wire_in_186 ),
       .io_V_wire_in_9( io_V_wire_in_185 ),
       .io_V_wire_in_8( io_V_wire_in_184 ),
       .io_V_wire_in_7( io_V_wire_in_183 ),
       .io_V_wire_in_6( io_V_wire_in_182 ),
       .io_V_wire_in_5( io_V_wire_in_181 ),
       .io_V_wire_in_4( io_V_wire_in_180 ),
       .io_V_wire_in_3( io_V_wire_in_179 ),
       .io_V_wire_in_2( io_V_wire_in_178 ),
       .io_V_wire_in_1( io_V_wire_in_177 ),
       .io_V_wire_in_0( io_V_wire_in_176 ),
       .io_H_wire_above_in_10( io_H_wire_above_21 ),
       .io_H_wire_above_in_9( io_H_wire_above_20 ),
       .io_H_wire_above_in_8( io_H_wire_above_19 ),
       .io_H_wire_above_in_7( io_H_wire_above_18 ),
       .io_H_wire_above_in_6( io_H_wire_above_17 ),
       .io_H_wire_above_in_5( io_H_wire_above_16 ),
       .io_H_wire_above_in_4( io_H_wire_above_15 ),
       .io_H_wire_above_in_3( io_H_wire_above_14 ),
       .io_H_wire_above_in_2( io_H_wire_above_13 ),
       .io_H_wire_above_in_1( io_H_wire_above_12 ),
       .io_H_wire_above_in_0( io_H_wire_above_11 ),
       .io_H_wire_below_in_10( H_wire_below_21 ),
       .io_H_wire_below_in_9( H_wire_below_20 ),
       .io_H_wire_below_in_8( H_wire_below_19 ),
       .io_H_wire_below_in_7( H_wire_below_18 ),
       .io_H_wire_below_in_6( H_wire_below_17 ),
       .io_H_wire_below_in_5( H_wire_below_16 ),
       .io_H_wire_below_in_4( H_wire_below_15 ),
       .io_H_wire_below_in_3( H_wire_below_14 ),
       .io_H_wire_below_in_2( H_wire_below_13 ),
       .io_H_wire_below_in_1( H_wire_below_12 ),
       .io_H_wire_below_in_0( H_wire_below_11 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_11 ),
       .io_shift_X_in_2( LogicBlockModule_10_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_10_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_10_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_11 ),
       .io_shift_carry_in( LogicBlockModule_10_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_10_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_11_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_11_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_11_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_11_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_11_io_carry_out ),
       .io_store_en( T1154 ),
       .io_mem_D_or_Z( T1149 ),
       .io_config( config_11 ),
       .io_mem_bus_out( LogicBlockModule_11_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_11_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_11_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_11_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_11_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_11_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_12(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_207 ),
       .io_V_wire_in_14( io_V_wire_in_206 ),
       .io_V_wire_in_13( io_V_wire_in_205 ),
       .io_V_wire_in_12( io_V_wire_in_204 ),
       .io_V_wire_in_11( io_V_wire_in_203 ),
       .io_V_wire_in_10( io_V_wire_in_202 ),
       .io_V_wire_in_9( io_V_wire_in_201 ),
       .io_V_wire_in_8( io_V_wire_in_200 ),
       .io_V_wire_in_7( io_V_wire_in_199 ),
       .io_V_wire_in_6( io_V_wire_in_198 ),
       .io_V_wire_in_5( io_V_wire_in_197 ),
       .io_V_wire_in_4( io_V_wire_in_196 ),
       .io_V_wire_in_3( io_V_wire_in_195 ),
       .io_V_wire_in_2( io_V_wire_in_194 ),
       .io_V_wire_in_1( io_V_wire_in_193 ),
       .io_V_wire_in_0( io_V_wire_in_192 ),
       .io_H_wire_above_in_10( io_H_wire_above_20 ),
       .io_H_wire_above_in_9( io_H_wire_above_19 ),
       .io_H_wire_above_in_8( io_H_wire_above_18 ),
       .io_H_wire_above_in_7( io_H_wire_above_17 ),
       .io_H_wire_above_in_6( io_H_wire_above_16 ),
       .io_H_wire_above_in_5( io_H_wire_above_15 ),
       .io_H_wire_above_in_4( io_H_wire_above_14 ),
       .io_H_wire_above_in_3( io_H_wire_above_13 ),
       .io_H_wire_above_in_2( io_H_wire_above_12 ),
       .io_H_wire_above_in_1( io_H_wire_above_11 ),
       .io_H_wire_above_in_0( io_H_wire_above_10 ),
       .io_H_wire_below_in_10( H_wire_below_20 ),
       .io_H_wire_below_in_9( H_wire_below_19 ),
       .io_H_wire_below_in_8( H_wire_below_18 ),
       .io_H_wire_below_in_7( H_wire_below_17 ),
       .io_H_wire_below_in_6( H_wire_below_16 ),
       .io_H_wire_below_in_5( H_wire_below_15 ),
       .io_H_wire_below_in_4( H_wire_below_14 ),
       .io_H_wire_below_in_3( H_wire_below_13 ),
       .io_H_wire_below_in_2( H_wire_below_12 ),
       .io_H_wire_below_in_1( H_wire_below_11 ),
       .io_H_wire_below_in_0( H_wire_below_10 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_12 ),
       .io_shift_X_in_2( LogicBlockModule_11_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_11_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_11_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_12 ),
       .io_shift_carry_in( LogicBlockModule_11_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_11_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_12_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_12_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_12_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_12_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_12_io_carry_out ),
       .io_store_en( T1146 ),
       .io_mem_D_or_Z( T1141 ),
       .io_config( config_12 ),
       .io_mem_bus_out( LogicBlockModule_12_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_12_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_12_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_12_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_12_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_12_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_13(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_223 ),
       .io_V_wire_in_14( io_V_wire_in_222 ),
       .io_V_wire_in_13( io_V_wire_in_221 ),
       .io_V_wire_in_12( io_V_wire_in_220 ),
       .io_V_wire_in_11( io_V_wire_in_219 ),
       .io_V_wire_in_10( io_V_wire_in_218 ),
       .io_V_wire_in_9( io_V_wire_in_217 ),
       .io_V_wire_in_8( io_V_wire_in_216 ),
       .io_V_wire_in_7( io_V_wire_in_215 ),
       .io_V_wire_in_6( io_V_wire_in_214 ),
       .io_V_wire_in_5( io_V_wire_in_213 ),
       .io_V_wire_in_4( io_V_wire_in_212 ),
       .io_V_wire_in_3( io_V_wire_in_211 ),
       .io_V_wire_in_2( io_V_wire_in_210 ),
       .io_V_wire_in_1( io_V_wire_in_209 ),
       .io_V_wire_in_0( io_V_wire_in_208 ),
       .io_H_wire_above_in_10( io_H_wire_above_19 ),
       .io_H_wire_above_in_9( io_H_wire_above_18 ),
       .io_H_wire_above_in_8( io_H_wire_above_17 ),
       .io_H_wire_above_in_7( io_H_wire_above_16 ),
       .io_H_wire_above_in_6( io_H_wire_above_15 ),
       .io_H_wire_above_in_5( io_H_wire_above_14 ),
       .io_H_wire_above_in_4( io_H_wire_above_13 ),
       .io_H_wire_above_in_3( io_H_wire_above_12 ),
       .io_H_wire_above_in_2( io_H_wire_above_11 ),
       .io_H_wire_above_in_1( io_H_wire_above_10 ),
       .io_H_wire_above_in_0( io_H_wire_above_9 ),
       .io_H_wire_below_in_10( H_wire_below_19 ),
       .io_H_wire_below_in_9( H_wire_below_18 ),
       .io_H_wire_below_in_8( H_wire_below_17 ),
       .io_H_wire_below_in_7( H_wire_below_16 ),
       .io_H_wire_below_in_6( H_wire_below_15 ),
       .io_H_wire_below_in_5( H_wire_below_14 ),
       .io_H_wire_below_in_4( H_wire_below_13 ),
       .io_H_wire_below_in_3( H_wire_below_12 ),
       .io_H_wire_below_in_2( H_wire_below_11 ),
       .io_H_wire_below_in_1( H_wire_below_10 ),
       .io_H_wire_below_in_0( H_wire_below_9 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_13 ),
       .io_shift_X_in_2( LogicBlockModule_12_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_12_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_12_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_13 ),
       .io_shift_carry_in( LogicBlockModule_12_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_12_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_13_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_13_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_13_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_13_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_13_io_carry_out ),
       .io_store_en( T1138 ),
       .io_mem_D_or_Z( T1133 ),
       .io_config( config_13 ),
       .io_mem_bus_out( LogicBlockModule_13_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_13_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_13_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_13_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_13_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_13_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_14(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_239 ),
       .io_V_wire_in_14( io_V_wire_in_238 ),
       .io_V_wire_in_13( io_V_wire_in_237 ),
       .io_V_wire_in_12( io_V_wire_in_236 ),
       .io_V_wire_in_11( io_V_wire_in_235 ),
       .io_V_wire_in_10( io_V_wire_in_234 ),
       .io_V_wire_in_9( io_V_wire_in_233 ),
       .io_V_wire_in_8( io_V_wire_in_232 ),
       .io_V_wire_in_7( io_V_wire_in_231 ),
       .io_V_wire_in_6( io_V_wire_in_230 ),
       .io_V_wire_in_5( io_V_wire_in_229 ),
       .io_V_wire_in_4( io_V_wire_in_228 ),
       .io_V_wire_in_3( io_V_wire_in_227 ),
       .io_V_wire_in_2( io_V_wire_in_226 ),
       .io_V_wire_in_1( io_V_wire_in_225 ),
       .io_V_wire_in_0( io_V_wire_in_224 ),
       .io_H_wire_above_in_10( io_H_wire_above_18 ),
       .io_H_wire_above_in_9( io_H_wire_above_17 ),
       .io_H_wire_above_in_8( io_H_wire_above_16 ),
       .io_H_wire_above_in_7( io_H_wire_above_15 ),
       .io_H_wire_above_in_6( io_H_wire_above_14 ),
       .io_H_wire_above_in_5( io_H_wire_above_13 ),
       .io_H_wire_above_in_4( io_H_wire_above_12 ),
       .io_H_wire_above_in_3( io_H_wire_above_11 ),
       .io_H_wire_above_in_2( io_H_wire_above_10 ),
       .io_H_wire_above_in_1( io_H_wire_above_9 ),
       .io_H_wire_above_in_0( io_H_wire_above_8 ),
       .io_H_wire_below_in_10( H_wire_below_18 ),
       .io_H_wire_below_in_9( H_wire_below_17 ),
       .io_H_wire_below_in_8( H_wire_below_16 ),
       .io_H_wire_below_in_7( H_wire_below_15 ),
       .io_H_wire_below_in_6( H_wire_below_14 ),
       .io_H_wire_below_in_5( H_wire_below_13 ),
       .io_H_wire_below_in_4( H_wire_below_12 ),
       .io_H_wire_below_in_3( H_wire_below_11 ),
       .io_H_wire_below_in_2( H_wire_below_10 ),
       .io_H_wire_below_in_1( H_wire_below_9 ),
       .io_H_wire_below_in_0( H_wire_below_8 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_14 ),
       .io_shift_X_in_2( LogicBlockModule_13_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_13_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_13_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_14 ),
       .io_shift_carry_in( LogicBlockModule_13_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_13_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_14_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_14_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_14_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_14_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_14_io_carry_out ),
       .io_store_en( T1130 ),
       .io_mem_D_or_Z( T1125 ),
       .io_config( config_14 ),
       .io_mem_bus_out( LogicBlockModule_14_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_14_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_14_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_14_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_14_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_14_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_15(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_255 ),
       .io_V_wire_in_14( io_V_wire_in_254 ),
       .io_V_wire_in_13( io_V_wire_in_253 ),
       .io_V_wire_in_12( io_V_wire_in_252 ),
       .io_V_wire_in_11( io_V_wire_in_251 ),
       .io_V_wire_in_10( io_V_wire_in_250 ),
       .io_V_wire_in_9( io_V_wire_in_249 ),
       .io_V_wire_in_8( io_V_wire_in_248 ),
       .io_V_wire_in_7( io_V_wire_in_247 ),
       .io_V_wire_in_6( io_V_wire_in_246 ),
       .io_V_wire_in_5( io_V_wire_in_245 ),
       .io_V_wire_in_4( io_V_wire_in_244 ),
       .io_V_wire_in_3( io_V_wire_in_243 ),
       .io_V_wire_in_2( io_V_wire_in_242 ),
       .io_V_wire_in_1( io_V_wire_in_241 ),
       .io_V_wire_in_0( io_V_wire_in_240 ),
       .io_H_wire_above_in_10( io_H_wire_above_17 ),
       .io_H_wire_above_in_9( io_H_wire_above_16 ),
       .io_H_wire_above_in_8( io_H_wire_above_15 ),
       .io_H_wire_above_in_7( io_H_wire_above_14 ),
       .io_H_wire_above_in_6( io_H_wire_above_13 ),
       .io_H_wire_above_in_5( io_H_wire_above_12 ),
       .io_H_wire_above_in_4( io_H_wire_above_11 ),
       .io_H_wire_above_in_3( io_H_wire_above_10 ),
       .io_H_wire_above_in_2( io_H_wire_above_9 ),
       .io_H_wire_above_in_1( io_H_wire_above_8 ),
       .io_H_wire_above_in_0( io_H_wire_above_7 ),
       .io_H_wire_below_in_10( H_wire_below_17 ),
       .io_H_wire_below_in_9( H_wire_below_16 ),
       .io_H_wire_below_in_8( H_wire_below_15 ),
       .io_H_wire_below_in_7( H_wire_below_14 ),
       .io_H_wire_below_in_6( H_wire_below_13 ),
       .io_H_wire_below_in_5( H_wire_below_12 ),
       .io_H_wire_below_in_4( H_wire_below_11 ),
       .io_H_wire_below_in_3( H_wire_below_10 ),
       .io_H_wire_below_in_2( H_wire_below_9 ),
       .io_H_wire_below_in_1( H_wire_below_8 ),
       .io_H_wire_below_in_0( H_wire_below_7 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_15 ),
       .io_shift_X_in_2( LogicBlockModule_14_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_14_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_14_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_15 ),
       .io_shift_carry_in( LogicBlockModule_14_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_14_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_15_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_15_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_15_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_15_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_15_io_carry_out ),
       .io_store_en( T1122 ),
       .io_mem_D_or_Z( T1117 ),
       .io_config( config_15 ),
       .io_mem_bus_out( LogicBlockModule_15_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_15_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_15_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_15_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_15_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_15_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_16(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_271 ),
       .io_V_wire_in_14( io_V_wire_in_270 ),
       .io_V_wire_in_13( io_V_wire_in_269 ),
       .io_V_wire_in_12( io_V_wire_in_268 ),
       .io_V_wire_in_11( io_V_wire_in_267 ),
       .io_V_wire_in_10( io_V_wire_in_266 ),
       .io_V_wire_in_9( io_V_wire_in_265 ),
       .io_V_wire_in_8( io_V_wire_in_264 ),
       .io_V_wire_in_7( io_V_wire_in_263 ),
       .io_V_wire_in_6( io_V_wire_in_262 ),
       .io_V_wire_in_5( io_V_wire_in_261 ),
       .io_V_wire_in_4( io_V_wire_in_260 ),
       .io_V_wire_in_3( io_V_wire_in_259 ),
       .io_V_wire_in_2( io_V_wire_in_258 ),
       .io_V_wire_in_1( io_V_wire_in_257 ),
       .io_V_wire_in_0( io_V_wire_in_256 ),
       .io_H_wire_above_in_10( io_H_wire_above_16 ),
       .io_H_wire_above_in_9( io_H_wire_above_15 ),
       .io_H_wire_above_in_8( io_H_wire_above_14 ),
       .io_H_wire_above_in_7( io_H_wire_above_13 ),
       .io_H_wire_above_in_6( io_H_wire_above_12 ),
       .io_H_wire_above_in_5( io_H_wire_above_11 ),
       .io_H_wire_above_in_4( io_H_wire_above_10 ),
       .io_H_wire_above_in_3( io_H_wire_above_9 ),
       .io_H_wire_above_in_2( io_H_wire_above_8 ),
       .io_H_wire_above_in_1( io_H_wire_above_7 ),
       .io_H_wire_above_in_0( io_H_wire_above_6 ),
       .io_H_wire_below_in_10( H_wire_below_16 ),
       .io_H_wire_below_in_9( H_wire_below_15 ),
       .io_H_wire_below_in_8( H_wire_below_14 ),
       .io_H_wire_below_in_7( H_wire_below_13 ),
       .io_H_wire_below_in_6( H_wire_below_12 ),
       .io_H_wire_below_in_5( H_wire_below_11 ),
       .io_H_wire_below_in_4( H_wire_below_10 ),
       .io_H_wire_below_in_3( H_wire_below_9 ),
       .io_H_wire_below_in_2( H_wire_below_8 ),
       .io_H_wire_below_in_1( H_wire_below_7 ),
       .io_H_wire_below_in_0( H_wire_below_6 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_16 ),
       .io_shift_X_in_2( LogicBlockModule_15_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_15_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_15_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_16 ),
       .io_shift_carry_in( LogicBlockModule_15_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_15_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_16_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_16_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_16_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_16_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_16_io_carry_out ),
       .io_store_en( T1114 ),
       .io_mem_D_or_Z( T1109 ),
       .io_config( config_16 ),
       .io_mem_bus_out( LogicBlockModule_16_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_16_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_16_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_16_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_16_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_16_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_17(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_287 ),
       .io_V_wire_in_14( io_V_wire_in_286 ),
       .io_V_wire_in_13( io_V_wire_in_285 ),
       .io_V_wire_in_12( io_V_wire_in_284 ),
       .io_V_wire_in_11( io_V_wire_in_283 ),
       .io_V_wire_in_10( io_V_wire_in_282 ),
       .io_V_wire_in_9( io_V_wire_in_281 ),
       .io_V_wire_in_8( io_V_wire_in_280 ),
       .io_V_wire_in_7( io_V_wire_in_279 ),
       .io_V_wire_in_6( io_V_wire_in_278 ),
       .io_V_wire_in_5( io_V_wire_in_277 ),
       .io_V_wire_in_4( io_V_wire_in_276 ),
       .io_V_wire_in_3( io_V_wire_in_275 ),
       .io_V_wire_in_2( io_V_wire_in_274 ),
       .io_V_wire_in_1( io_V_wire_in_273 ),
       .io_V_wire_in_0( io_V_wire_in_272 ),
       .io_H_wire_above_in_10( io_H_wire_above_15 ),
       .io_H_wire_above_in_9( io_H_wire_above_14 ),
       .io_H_wire_above_in_8( io_H_wire_above_13 ),
       .io_H_wire_above_in_7( io_H_wire_above_12 ),
       .io_H_wire_above_in_6( io_H_wire_above_11 ),
       .io_H_wire_above_in_5( io_H_wire_above_10 ),
       .io_H_wire_above_in_4( io_H_wire_above_9 ),
       .io_H_wire_above_in_3( io_H_wire_above_8 ),
       .io_H_wire_above_in_2( io_H_wire_above_7 ),
       .io_H_wire_above_in_1( io_H_wire_above_6 ),
       .io_H_wire_above_in_0( io_H_wire_above_5 ),
       .io_H_wire_below_in_10( H_wire_below_15 ),
       .io_H_wire_below_in_9( H_wire_below_14 ),
       .io_H_wire_below_in_8( H_wire_below_13 ),
       .io_H_wire_below_in_7( H_wire_below_12 ),
       .io_H_wire_below_in_6( H_wire_below_11 ),
       .io_H_wire_below_in_5( H_wire_below_10 ),
       .io_H_wire_below_in_4( H_wire_below_9 ),
       .io_H_wire_below_in_3( H_wire_below_8 ),
       .io_H_wire_below_in_2( H_wire_below_7 ),
       .io_H_wire_below_in_1( H_wire_below_6 ),
       .io_H_wire_below_in_0( H_wire_below_5 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_17 ),
       .io_shift_X_in_2( LogicBlockModule_16_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_16_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_16_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_17 ),
       .io_shift_carry_in( LogicBlockModule_16_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_16_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_17_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_17_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_17_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_17_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_17_io_carry_out ),
       .io_store_en( T1106 ),
       .io_mem_D_or_Z( T1101 ),
       .io_config( config_17 ),
       .io_mem_bus_out( LogicBlockModule_17_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_17_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_17_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_17_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_17_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_17_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_18(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_303 ),
       .io_V_wire_in_14( io_V_wire_in_302 ),
       .io_V_wire_in_13( io_V_wire_in_301 ),
       .io_V_wire_in_12( io_V_wire_in_300 ),
       .io_V_wire_in_11( io_V_wire_in_299 ),
       .io_V_wire_in_10( io_V_wire_in_298 ),
       .io_V_wire_in_9( io_V_wire_in_297 ),
       .io_V_wire_in_8( io_V_wire_in_296 ),
       .io_V_wire_in_7( io_V_wire_in_295 ),
       .io_V_wire_in_6( io_V_wire_in_294 ),
       .io_V_wire_in_5( io_V_wire_in_293 ),
       .io_V_wire_in_4( io_V_wire_in_292 ),
       .io_V_wire_in_3( io_V_wire_in_291 ),
       .io_V_wire_in_2( io_V_wire_in_290 ),
       .io_V_wire_in_1( io_V_wire_in_289 ),
       .io_V_wire_in_0( io_V_wire_in_288 ),
       .io_H_wire_above_in_10( io_H_wire_above_14 ),
       .io_H_wire_above_in_9( io_H_wire_above_13 ),
       .io_H_wire_above_in_8( io_H_wire_above_12 ),
       .io_H_wire_above_in_7( io_H_wire_above_11 ),
       .io_H_wire_above_in_6( io_H_wire_above_10 ),
       .io_H_wire_above_in_5( io_H_wire_above_9 ),
       .io_H_wire_above_in_4( io_H_wire_above_8 ),
       .io_H_wire_above_in_3( io_H_wire_above_7 ),
       .io_H_wire_above_in_2( io_H_wire_above_6 ),
       .io_H_wire_above_in_1( io_H_wire_above_5 ),
       .io_H_wire_above_in_0( io_H_wire_above_4 ),
       .io_H_wire_below_in_10( H_wire_below_14 ),
       .io_H_wire_below_in_9( H_wire_below_13 ),
       .io_H_wire_below_in_8( H_wire_below_12 ),
       .io_H_wire_below_in_7( H_wire_below_11 ),
       .io_H_wire_below_in_6( H_wire_below_10 ),
       .io_H_wire_below_in_5( H_wire_below_9 ),
       .io_H_wire_below_in_4( H_wire_below_8 ),
       .io_H_wire_below_in_3( H_wire_below_7 ),
       .io_H_wire_below_in_2( H_wire_below_6 ),
       .io_H_wire_below_in_1( H_wire_below_5 ),
       .io_H_wire_below_in_0( H_wire_below_4 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_18 ),
       .io_shift_X_in_2( LogicBlockModule_17_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_17_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_17_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_18 ),
       .io_shift_carry_in( LogicBlockModule_17_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_17_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_18_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_18_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_18_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_18_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_18_io_carry_out ),
       .io_store_en( T1098 ),
       .io_mem_D_or_Z( T1093 ),
       .io_config( config_18 ),
       .io_mem_bus_out( LogicBlockModule_18_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_18_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_18_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_18_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_18_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_18_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_19(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_319 ),
       .io_V_wire_in_14( io_V_wire_in_318 ),
       .io_V_wire_in_13( io_V_wire_in_317 ),
       .io_V_wire_in_12( io_V_wire_in_316 ),
       .io_V_wire_in_11( io_V_wire_in_315 ),
       .io_V_wire_in_10( io_V_wire_in_314 ),
       .io_V_wire_in_9( io_V_wire_in_313 ),
       .io_V_wire_in_8( io_V_wire_in_312 ),
       .io_V_wire_in_7( io_V_wire_in_311 ),
       .io_V_wire_in_6( io_V_wire_in_310 ),
       .io_V_wire_in_5( io_V_wire_in_309 ),
       .io_V_wire_in_4( io_V_wire_in_308 ),
       .io_V_wire_in_3( io_V_wire_in_307 ),
       .io_V_wire_in_2( io_V_wire_in_306 ),
       .io_V_wire_in_1( io_V_wire_in_305 ),
       .io_V_wire_in_0( io_V_wire_in_304 ),
       .io_H_wire_above_in_10( io_H_wire_above_13 ),
       .io_H_wire_above_in_9( io_H_wire_above_12 ),
       .io_H_wire_above_in_8( io_H_wire_above_11 ),
       .io_H_wire_above_in_7( io_H_wire_above_10 ),
       .io_H_wire_above_in_6( io_H_wire_above_9 ),
       .io_H_wire_above_in_5( io_H_wire_above_8 ),
       .io_H_wire_above_in_4( io_H_wire_above_7 ),
       .io_H_wire_above_in_3( io_H_wire_above_6 ),
       .io_H_wire_above_in_2( io_H_wire_above_5 ),
       .io_H_wire_above_in_1( io_H_wire_above_4 ),
       .io_H_wire_above_in_0( io_H_wire_above_3 ),
       .io_H_wire_below_in_10( H_wire_below_13 ),
       .io_H_wire_below_in_9( H_wire_below_12 ),
       .io_H_wire_below_in_8( H_wire_below_11 ),
       .io_H_wire_below_in_7( H_wire_below_10 ),
       .io_H_wire_below_in_6( H_wire_below_9 ),
       .io_H_wire_below_in_5( H_wire_below_8 ),
       .io_H_wire_below_in_4( H_wire_below_7 ),
       .io_H_wire_below_in_3( H_wire_below_6 ),
       .io_H_wire_below_in_2( H_wire_below_5 ),
       .io_H_wire_below_in_1( H_wire_below_4 ),
       .io_H_wire_below_in_0( H_wire_below_3 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_19 ),
       .io_shift_X_in_2( LogicBlockModule_18_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_18_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_18_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_19 ),
       .io_shift_carry_in( LogicBlockModule_18_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_18_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_19_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_19_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_19_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_19_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_19_io_carry_out ),
       .io_store_en( T1090 ),
       .io_mem_D_or_Z( T1085 ),
       .io_config( config_19 ),
       .io_mem_bus_out( LogicBlockModule_19_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_19_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_19_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_19_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_19_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_19_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_20(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_335 ),
       .io_V_wire_in_14( io_V_wire_in_334 ),
       .io_V_wire_in_13( io_V_wire_in_333 ),
       .io_V_wire_in_12( io_V_wire_in_332 ),
       .io_V_wire_in_11( io_V_wire_in_331 ),
       .io_V_wire_in_10( io_V_wire_in_330 ),
       .io_V_wire_in_9( io_V_wire_in_329 ),
       .io_V_wire_in_8( io_V_wire_in_328 ),
       .io_V_wire_in_7( io_V_wire_in_327 ),
       .io_V_wire_in_6( io_V_wire_in_326 ),
       .io_V_wire_in_5( io_V_wire_in_325 ),
       .io_V_wire_in_4( io_V_wire_in_324 ),
       .io_V_wire_in_3( io_V_wire_in_323 ),
       .io_V_wire_in_2( io_V_wire_in_322 ),
       .io_V_wire_in_1( io_V_wire_in_321 ),
       .io_V_wire_in_0( io_V_wire_in_320 ),
       .io_H_wire_above_in_10( io_H_wire_above_12 ),
       .io_H_wire_above_in_9( io_H_wire_above_11 ),
       .io_H_wire_above_in_8( io_H_wire_above_10 ),
       .io_H_wire_above_in_7( io_H_wire_above_9 ),
       .io_H_wire_above_in_6( io_H_wire_above_8 ),
       .io_H_wire_above_in_5( io_H_wire_above_7 ),
       .io_H_wire_above_in_4( io_H_wire_above_6 ),
       .io_H_wire_above_in_3( io_H_wire_above_5 ),
       .io_H_wire_above_in_2( io_H_wire_above_4 ),
       .io_H_wire_above_in_1( io_H_wire_above_3 ),
       .io_H_wire_above_in_0( io_H_wire_above_2 ),
       .io_H_wire_below_in_10( H_wire_below_12 ),
       .io_H_wire_below_in_9( H_wire_below_11 ),
       .io_H_wire_below_in_8( H_wire_below_10 ),
       .io_H_wire_below_in_7( H_wire_below_9 ),
       .io_H_wire_below_in_6( H_wire_below_8 ),
       .io_H_wire_below_in_5( H_wire_below_7 ),
       .io_H_wire_below_in_4( H_wire_below_6 ),
       .io_H_wire_below_in_3( H_wire_below_5 ),
       .io_H_wire_below_in_2( H_wire_below_4 ),
       .io_H_wire_below_in_1( H_wire_below_3 ),
       .io_H_wire_below_in_0( H_wire_below_2 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_20 ),
       .io_shift_X_in_2( LogicBlockModule_19_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_19_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_19_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_20 ),
       .io_shift_carry_in( LogicBlockModule_19_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_19_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_20_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_20_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_20_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_20_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_20_io_carry_out ),
       .io_store_en( T1082 ),
       .io_mem_D_or_Z( T1077 ),
       .io_config( config_20 ),
       .io_mem_bus_out( LogicBlockModule_20_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_20_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_20_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_20_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_20_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_20_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_21(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_351 ),
       .io_V_wire_in_14( io_V_wire_in_350 ),
       .io_V_wire_in_13( io_V_wire_in_349 ),
       .io_V_wire_in_12( io_V_wire_in_348 ),
       .io_V_wire_in_11( io_V_wire_in_347 ),
       .io_V_wire_in_10( io_V_wire_in_346 ),
       .io_V_wire_in_9( io_V_wire_in_345 ),
       .io_V_wire_in_8( io_V_wire_in_344 ),
       .io_V_wire_in_7( io_V_wire_in_343 ),
       .io_V_wire_in_6( io_V_wire_in_342 ),
       .io_V_wire_in_5( io_V_wire_in_341 ),
       .io_V_wire_in_4( io_V_wire_in_340 ),
       .io_V_wire_in_3( io_V_wire_in_339 ),
       .io_V_wire_in_2( io_V_wire_in_338 ),
       .io_V_wire_in_1( io_V_wire_in_337 ),
       .io_V_wire_in_0( io_V_wire_in_336 ),
       .io_H_wire_above_in_10( io_H_wire_above_11 ),
       .io_H_wire_above_in_9( io_H_wire_above_10 ),
       .io_H_wire_above_in_8( io_H_wire_above_9 ),
       .io_H_wire_above_in_7( io_H_wire_above_8 ),
       .io_H_wire_above_in_6( io_H_wire_above_7 ),
       .io_H_wire_above_in_5( io_H_wire_above_6 ),
       .io_H_wire_above_in_4( io_H_wire_above_5 ),
       .io_H_wire_above_in_3( io_H_wire_above_4 ),
       .io_H_wire_above_in_2( io_H_wire_above_3 ),
       .io_H_wire_above_in_1( io_H_wire_above_2 ),
       .io_H_wire_above_in_0( io_H_wire_above_1 ),
       .io_H_wire_below_in_10( H_wire_below_11 ),
       .io_H_wire_below_in_9( H_wire_below_10 ),
       .io_H_wire_below_in_8( H_wire_below_9 ),
       .io_H_wire_below_in_7( H_wire_below_8 ),
       .io_H_wire_below_in_6( H_wire_below_7 ),
       .io_H_wire_below_in_5( H_wire_below_6 ),
       .io_H_wire_below_in_4( H_wire_below_5 ),
       .io_H_wire_below_in_3( H_wire_below_4 ),
       .io_H_wire_below_in_2( H_wire_below_3 ),
       .io_H_wire_below_in_1( H_wire_below_2 ),
       .io_H_wire_below_in_0( H_wire_below_1 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_21 ),
       .io_shift_X_in_2( LogicBlockModule_20_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_20_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_20_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_21 ),
       .io_shift_carry_in( LogicBlockModule_20_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_20_io_carry_out ),
       .io_shift_X_out_2( LogicBlockModule_21_io_shift_X_out_2 ),
       .io_shift_X_out_1( LogicBlockModule_21_io_shift_X_out_1 ),
       .io_shift_X_out_0( LogicBlockModule_21_io_shift_X_out_0 ),
       .io_shift_carry_out( LogicBlockModule_21_io_shift_carry_out ),
       .io_carry_out( LogicBlockModule_21_io_carry_out ),
       .io_store_en( T1074 ),
       .io_mem_D_or_Z( T1069 ),
       .io_config( config_21 ),
       .io_mem_bus_out( LogicBlockModule_21_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_21_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_21_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_21_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_21_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_21_io_config_V_out )
  );
  LogicBlockModule LogicBlockModule_22(.clk(clk), .reset(reset),
       .io_V_wire_in_15( io_V_wire_in_367 ),
       .io_V_wire_in_14( io_V_wire_in_366 ),
       .io_V_wire_in_13( io_V_wire_in_365 ),
       .io_V_wire_in_12( io_V_wire_in_364 ),
       .io_V_wire_in_11( io_V_wire_in_363 ),
       .io_V_wire_in_10( io_V_wire_in_362 ),
       .io_V_wire_in_9( io_V_wire_in_361 ),
       .io_V_wire_in_8( io_V_wire_in_360 ),
       .io_V_wire_in_7( io_V_wire_in_359 ),
       .io_V_wire_in_6( io_V_wire_in_358 ),
       .io_V_wire_in_5( io_V_wire_in_357 ),
       .io_V_wire_in_4( io_V_wire_in_356 ),
       .io_V_wire_in_3( io_V_wire_in_355 ),
       .io_V_wire_in_2( io_V_wire_in_354 ),
       .io_V_wire_in_1( io_V_wire_in_353 ),
       .io_V_wire_in_0( io_V_wire_in_352 ),
       .io_H_wire_above_in_10( io_H_wire_above_10 ),
       .io_H_wire_above_in_9( io_H_wire_above_9 ),
       .io_H_wire_above_in_8( io_H_wire_above_8 ),
       .io_H_wire_above_in_7( io_H_wire_above_7 ),
       .io_H_wire_above_in_6( io_H_wire_above_6 ),
       .io_H_wire_above_in_5( io_H_wire_above_5 ),
       .io_H_wire_above_in_4( io_H_wire_above_4 ),
       .io_H_wire_above_in_3( io_H_wire_above_3 ),
       .io_H_wire_above_in_2( io_H_wire_above_2 ),
       .io_H_wire_above_in_1( io_H_wire_above_1 ),
       .io_H_wire_above_in_0( io_H_wire_above_0 ),
       .io_H_wire_below_in_10( H_wire_below_10 ),
       .io_H_wire_below_in_9( H_wire_below_9 ),
       .io_H_wire_below_in_8( H_wire_below_8 ),
       .io_H_wire_below_in_7( H_wire_below_7 ),
       .io_H_wire_below_in_6( H_wire_below_6 ),
       .io_H_wire_below_in_5( H_wire_below_5 ),
       .io_H_wire_below_in_4( H_wire_below_4 ),
       .io_H_wire_below_in_3( H_wire_below_3 ),
       .io_H_wire_below_in_2( H_wire_below_2 ),
       .io_H_wire_below_in_1( H_wire_below_1 ),
       .io_H_wire_below_in_0( H_wire_below_0 ),
       .io_G_wire_above_in_3( io_G_wire_above_3 ),
       .io_G_wire_above_in_2( io_G_wire_above_2 ),
       .io_G_wire_above_in_1( io_G_wire_above_1 ),
       .io_G_wire_above_in_0( io_G_wire_above_0 ),
       .io_G_wire_below_in_3( G_wire_below_3 ),
       .io_G_wire_below_in_2( G_wire_below_2 ),
       .io_G_wire_below_in_1( G_wire_below_1 ),
       .io_G_wire_below_in_0( G_wire_below_0 ),
       .io_mem_bus_in( io_mem_bus_in_22 ),
       .io_shift_X_in_2( LogicBlockModule_21_io_shift_X_out_2 ),
       .io_shift_X_in_1( LogicBlockModule_21_io_shift_X_out_1 ),
       .io_shift_X_in_0( LogicBlockModule_21_io_shift_X_out_0 ),
       .io_H_out_above( io_H_out_above_22 ),
       .io_shift_carry_in( LogicBlockModule_21_io_shift_carry_out ),
       .io_carry_in( LogicBlockModule_21_io_carry_out ),
       //.io_shift_X_out_2(  )
       //.io_shift_X_out_1(  )
       //.io_shift_X_out_0(  )
       //.io_shift_carry_out(  )
       //.io_carry_out(  )
       .io_store_en( T1066 ),
       .io_mem_D_or_Z( T1061 ),
       .io_config( config_22 ),
       .io_mem_bus_out( LogicBlockModule_22_io_mem_bus_out ),
       .io_V_wire_out( LogicBlockModule_22_io_V_wire_out ),
       .io_H_wire_out( LogicBlockModule_22_io_H_wire_out ),
       .io_G_wire_out( LogicBlockModule_22_io_G_wire_out ),
       .io_config_G_out( LogicBlockModule_22_io_config_G_out ),
       .io_config_V_out( LogicBlockModule_22_io_config_V_out )
  );
  GWireModule GWireModule(
       .io_G_in_22( G_wire_outs_22 ),
       .io_G_in_21( G_wire_outs_21 ),
       .io_G_in_20( G_wire_outs_20 ),
       .io_G_in_19( G_wire_outs_19 ),
       .io_G_in_18( G_wire_outs_18 ),
       .io_G_in_17( G_wire_outs_17 ),
       .io_G_in_16( G_wire_outs_16 ),
       .io_G_in_15( G_wire_outs_15 ),
       .io_G_in_14( G_wire_outs_14 ),
       .io_G_in_13( G_wire_outs_13 ),
       .io_G_in_12( G_wire_outs_12 ),
       .io_G_in_11( G_wire_outs_11 ),
       .io_G_in_10( G_wire_outs_10 ),
       .io_G_in_9( G_wire_outs_9 ),
       .io_G_in_8( G_wire_outs_8 ),
       .io_G_in_7( G_wire_outs_7 ),
       .io_G_in_6( G_wire_outs_6 ),
       .io_G_in_5( G_wire_outs_5 ),
       .io_G_in_4( G_wire_outs_4 ),
       .io_G_in_3( G_wire_outs_3 ),
       .io_G_in_2( G_wire_outs_2 ),
       .io_G_in_1( G_wire_outs_1 ),
       .io_G_in_0( G_wire_outs_0 ),
       .io_en( G_wire_below_en_0 ),
       .io_G_out( GWireModule_io_G_out )
  );
  GWireModule GWireModule_1(
       .io_G_in_22( G_wire_outs_22 ),
       .io_G_in_21( G_wire_outs_21 ),
       .io_G_in_20( G_wire_outs_20 ),
       .io_G_in_19( G_wire_outs_19 ),
       .io_G_in_18( G_wire_outs_18 ),
       .io_G_in_17( G_wire_outs_17 ),
       .io_G_in_16( G_wire_outs_16 ),
       .io_G_in_15( G_wire_outs_15 ),
       .io_G_in_14( G_wire_outs_14 ),
       .io_G_in_13( G_wire_outs_13 ),
       .io_G_in_12( G_wire_outs_12 ),
       .io_G_in_11( G_wire_outs_11 ),
       .io_G_in_10( G_wire_outs_10 ),
       .io_G_in_9( G_wire_outs_9 ),
       .io_G_in_8( G_wire_outs_8 ),
       .io_G_in_7( G_wire_outs_7 ),
       .io_G_in_6( G_wire_outs_6 ),
       .io_G_in_5( G_wire_outs_5 ),
       .io_G_in_4( G_wire_outs_4 ),
       .io_G_in_3( G_wire_outs_3 ),
       .io_G_in_2( G_wire_outs_2 ),
       .io_G_in_1( G_wire_outs_1 ),
       .io_G_in_0( G_wire_outs_0 ),
       .io_en( G_wire_below_en_1 ),
       .io_G_out( GWireModule_1_io_G_out )
  );
  GWireModule GWireModule_2(
       .io_G_in_22( G_wire_outs_22 ),
       .io_G_in_21( G_wire_outs_21 ),
       .io_G_in_20( G_wire_outs_20 ),
       .io_G_in_19( G_wire_outs_19 ),
       .io_G_in_18( G_wire_outs_18 ),
       .io_G_in_17( G_wire_outs_17 ),
       .io_G_in_16( G_wire_outs_16 ),
       .io_G_in_15( G_wire_outs_15 ),
       .io_G_in_14( G_wire_outs_14 ),
       .io_G_in_13( G_wire_outs_13 ),
       .io_G_in_12( G_wire_outs_12 ),
       .io_G_in_11( G_wire_outs_11 ),
       .io_G_in_10( G_wire_outs_10 ),
       .io_G_in_9( G_wire_outs_9 ),
       .io_G_in_8( G_wire_outs_8 ),
       .io_G_in_7( G_wire_outs_7 ),
       .io_G_in_6( G_wire_outs_6 ),
       .io_G_in_5( G_wire_outs_5 ),
       .io_G_in_4( G_wire_outs_4 ),
       .io_G_in_3( G_wire_outs_3 ),
       .io_G_in_2( G_wire_outs_2 ),
       .io_G_in_1( G_wire_outs_1 ),
       .io_G_in_0( G_wire_outs_0 ),
       .io_en( G_wire_below_en_2 ),
       .io_G_out( GWireModule_2_io_G_out )
  );
  GWireModule GWireModule_3(
       .io_G_in_22( G_wire_outs_22 ),
       .io_G_in_21( G_wire_outs_21 ),
       .io_G_in_20( G_wire_outs_20 ),
       .io_G_in_19( G_wire_outs_19 ),
       .io_G_in_18( G_wire_outs_18 ),
       .io_G_in_17( G_wire_outs_17 ),
       .io_G_in_16( G_wire_outs_16 ),
       .io_G_in_15( G_wire_outs_15 ),
       .io_G_in_14( G_wire_outs_14 ),
       .io_G_in_13( G_wire_outs_13 ),
       .io_G_in_12( G_wire_outs_12 ),
       .io_G_in_11( G_wire_outs_11 ),
       .io_G_in_10( G_wire_outs_10 ),
       .io_G_in_9( G_wire_outs_9 ),
       .io_G_in_8( G_wire_outs_8 ),
       .io_G_in_7( G_wire_outs_7 ),
       .io_G_in_6( G_wire_outs_6 ),
       .io_G_in_5( G_wire_outs_5 ),
       .io_G_in_4( G_wire_outs_4 ),
       .io_G_in_3( G_wire_outs_3 ),
       .io_G_in_2( G_wire_outs_2 ),
       .io_G_in_1( G_wire_outs_1 ),
       .io_G_in_0( G_wire_outs_0 ),
       .io_en( G_wire_below_en_3 ),
       .io_G_out( GWireModule_3_io_G_out )
  );
  loop_wire LoopWireBlackBox(
       .in( GWireModule_io_G_out ),
       .out( LoopWireBlackBox_out )
  );
  loop_wire LoopWireBlackBox_1(
       .in( GWireModule_1_io_G_out ),
       .out( LoopWireBlackBox_1_out )
  );
  loop_wire LoopWireBlackBox_2(
       .in( GWireModule_2_io_G_out ),
       .out( LoopWireBlackBox_2_out )
  );
  loop_wire LoopWireBlackBox_3(
       .in( GWireModule_3_io_G_out ),
       .out( LoopWireBlackBox_3_out )
  );
  loop_wire LoopWireBlackBox_4(
       .in( 2'h0 ),
       .out( LoopWireBlackBox_4_out )
  );
  loop_wire LoopWireBlackBox_5(
       .in( T71 ),
       .out( LoopWireBlackBox_5_out )
  );
  loop_wire LoopWireBlackBox_6(
       .in( T70 ),
       .out( LoopWireBlackBox_6_out )
  );
  loop_wire LoopWireBlackBox_7(
       .in( T69 ),
       .out( LoopWireBlackBox_7_out )
  );
  loop_wire LoopWireBlackBox_8(
       .in( T68 ),
       .out( LoopWireBlackBox_8_out )
  );
  loop_wire LoopWireBlackBox_9(
       .in( T66 ),
       .out( LoopWireBlackBox_9_out )
  );
  loop_wire LoopWireBlackBox_10(
       .in( T64 ),
       .out( LoopWireBlackBox_10_out )
  );
  loop_wire LoopWireBlackBox_11(
       .in( T62 ),
       .out( LoopWireBlackBox_11_out )
  );
  loop_wire LoopWireBlackBox_12(
       .in( T60 ),
       .out( LoopWireBlackBox_12_out )
  );
  loop_wire LoopWireBlackBox_13(
       .in( T57 ),
       .out( LoopWireBlackBox_13_out )
  );
  loop_wire LoopWireBlackBox_14(
       .in( T54 ),
       .out( LoopWireBlackBox_14_out )
  );
  loop_wire LoopWireBlackBox_15(
       .in( T51 ),
       .out( LoopWireBlackBox_15_out )
  );
  loop_wire LoopWireBlackBox_16(
       .in( T48 ),
       .out( LoopWireBlackBox_16_out )
  );
  loop_wire LoopWireBlackBox_17(
       .in( T45 ),
       .out( LoopWireBlackBox_17_out )
  );
  loop_wire LoopWireBlackBox_18(
       .in( T42 ),
       .out( LoopWireBlackBox_18_out )
  );
  loop_wire LoopWireBlackBox_19(
       .in( T39 ),
       .out( LoopWireBlackBox_19_out )
  );
  loop_wire LoopWireBlackBox_20(
       .in( T36 ),
       .out( LoopWireBlackBox_20_out )
  );
  loop_wire LoopWireBlackBox_21(
       .in( T33 ),
       .out( LoopWireBlackBox_21_out )
  );
  loop_wire LoopWireBlackBox_22(
       .in( T30 ),
       .out( LoopWireBlackBox_22_out )
  );
  loop_wire LoopWireBlackBox_23(
       .in( T27 ),
       .out( LoopWireBlackBox_23_out )
  );
  loop_wire LoopWireBlackBox_24(
       .in( T24 ),
       .out( LoopWireBlackBox_24_out )
  );
  loop_wire LoopWireBlackBox_25(
       .in( T21 ),
       .out( LoopWireBlackBox_25_out )
  );
  loop_wire LoopWireBlackBox_26(
       .in( T18 ),
       .out( LoopWireBlackBox_26_out )
  );
  loop_wire LoopWireBlackBox_27(
       .in( T14 ),
       .out( LoopWireBlackBox_27_out )
  );
  loop_wire LoopWireBlackBox_28(
       .in( T12 ),
       .out( LoopWireBlackBox_28_out )
  );
  loop_wire LoopWireBlackBox_29(
       .in( T10 ),
       .out( LoopWireBlackBox_29_out )
  );
  loop_wire LoopWireBlackBox_30(
       .in( T8 ),
       .out( LoopWireBlackBox_30_out )
  );
  loop_wire LoopWireBlackBox_31(
       .in( T5 ),
       .out( LoopWireBlackBox_31_out )
  );
  loop_wire LoopWireBlackBox_32(
       .in( T4 ),
       .out( LoopWireBlackBox_32_out )
  );
  loop_wire LoopWireBlackBox_33(
       .in( T3 ),
       .out( LoopWireBlackBox_33_out )
  );
  loop_wire LoopWireBlackBox_34(
       .in( T2 ),
       .out( LoopWireBlackBox_34_out )
  );
  loop_wire LoopWireBlackBox_35(
       .in( T0 ),
       .out( LoopWireBlackBox_35_out )
  );
  loop_wire LoopWireBlackBox_36(
       .in( 2'h0 ),
       .out( LoopWireBlackBox_36_out )
  );
endmodule

module VwireBlackBox_0(
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    input  io_en_1,
    input  io_en_0,
    output[1:0] io_out
);

  wire[1:0] T26;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T27;
  wire T3;
  wire T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T28;
  wire[1:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T29;
  wire T10;
  wire T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[3:0] T30;
  wire[4:0] T14;
  wire[4:0] T31;
  wire[3:0] T15;
  wire[1:0] T16;
  wire[4:0] T17;
  wire[4:0] T18;
  wire[4:0] T19;
  wire[4:0] T32;
  wire[2:0] T20;
  wire[2:0] T33;
  wire[1:0] T21;
  wire[1:0] T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[1:0] VwireFlatBlackBox_out;


  assign T26 = T0[1'h1:1'h0];
  assign T0 = T5 | T1;
  assign T1 = T27 & T2;
  assign T2 = 3'h2;
  assign T27 = T3 ? 3'h7 : 3'h0;
  assign T3 = T4;
  assign T4 = io_en_1;
  assign T5 = T28 & T6;
  assign T6 = ~ T2;
  assign T28 = {1'h0, T7};
  assign T7 = T12 | T8;
  assign T8 = T29 & T9;
  assign T9 = 2'h1;
  assign T29 = T10 ? 2'h3 : 2'h0;
  assign T10 = T11;
  assign T11 = io_en_0;
  assign T12 = 2'h0 & T13;
  assign T13 = ~ T9;
  assign T30 = T14[2'h3:1'h0];
  assign T14 = T17 | T31;
  assign T31 = {1'h0, T15};
  assign T15 = T16 << 2'h2;
  assign T16 = io_in_1 & 2'h3;
  assign T17 = T32 & T18;
  assign T18 = ~ T19;
  assign T19 = 5'hc;
  assign T32 = {2'h0, T20};
  assign T20 = T23 | T33;
  assign T33 = {1'h0, T21};
  assign T21 = T22 << 1'h0;
  assign T22 = io_in_0 & 2'h3;
  assign T23 = 3'h0 & T24;
  assign T24 = ~ T25;
  assign T25 = 3'h3;
  assign io_out = VwireFlatBlackBox_out;
  vwire #(.W(2),.L(2)) VwireFlatBlackBox(
       .in( T30 ),
       .en( T26 ),
       .out( VwireFlatBlackBox_out )
  );
endmodule

module Vwire2BB(
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    input  io_en_1,
    input  io_en_0,
    output[1:0] io_out
);

  wire[1:0] VwireBlackBox_io_out;


  assign io_out = VwireBlackBox_io_out;
  VwireBlackBox_0 VwireBlackBox(
       .io_in_1( io_in_1 ),
       .io_in_0( io_in_0 ),
       .io_en_1( io_en_1 ),
       .io_en_0( io_en_0 ),
       .io_out( VwireBlackBox_io_out )
  );
endmodule

module Vwire_0(
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    input  io_en_1,
    input  io_en_0,
    output[1:0] io_out
);

  wire[1:0] Vwire2BB_io_out;


  assign io_out = Vwire2BB_io_out;
  Vwire2BB Vwire2BB(
       .io_in_1( io_in_1 ),
       .io_in_0( io_in_0 ),
       .io_en_1( io_en_1 ),
       .io_en_0( io_en_0 ),
       .io_out( Vwire2BB_io_out )
  );
endmodule

module VwireBlackBox_1(
    input [1:0] io_in_2,
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    input  io_en_2,
    input  io_en_1,
    input  io_en_0,
    output[1:0] io_out
);

  wire[2:0] T39;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T40;
  wire T3;
  wire T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T41;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T42;
  wire T10;
  wire T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T43;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire[1:0] T44;
  wire T17;
  wire T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[5:0] T45;
  wire[6:0] T21;
  wire[6:0] T46;
  wire[5:0] T22;
  wire[1:0] T23;
  wire[6:0] T24;
  wire[6:0] T25;
  wire[6:0] T26;
  wire[6:0] T47;
  wire[4:0] T27;
  wire[4:0] T48;
  wire[3:0] T28;
  wire[1:0] T29;
  wire[4:0] T30;
  wire[4:0] T31;
  wire[4:0] T32;
  wire[4:0] T49;
  wire[2:0] T33;
  wire[2:0] T50;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire[2:0] T38;
  wire[1:0] VwireFlatBlackBox_out;


  assign T39 = T0[2'h2:1'h0];
  assign T0 = T5 | T1;
  assign T1 = T40 & T2;
  assign T2 = 4'h4;
  assign T40 = T3 ? 4'hf : 4'h0;
  assign T3 = T4;
  assign T4 = io_en_2;
  assign T5 = T41 & T6;
  assign T6 = ~ T2;
  assign T41 = {1'h0, T7};
  assign T7 = T12 | T8;
  assign T8 = T42 & T9;
  assign T9 = 3'h2;
  assign T42 = T10 ? 3'h7 : 3'h0;
  assign T10 = T11;
  assign T11 = io_en_1;
  assign T12 = T43 & T13;
  assign T13 = ~ T9;
  assign T43 = {1'h0, T14};
  assign T14 = T19 | T15;
  assign T15 = T44 & T16;
  assign T16 = 2'h1;
  assign T44 = T17 ? 2'h3 : 2'h0;
  assign T17 = T18;
  assign T18 = io_en_0;
  assign T19 = 2'h0 & T20;
  assign T20 = ~ T16;
  assign T45 = T21[3'h5:1'h0];
  assign T21 = T24 | T46;
  assign T46 = {1'h0, T22};
  assign T22 = T23 << 3'h4;
  assign T23 = io_in_2 & 2'h3;
  assign T24 = T47 & T25;
  assign T25 = ~ T26;
  assign T26 = 7'h30;
  assign T47 = {2'h0, T27};
  assign T27 = T30 | T48;
  assign T48 = {1'h0, T28};
  assign T28 = T29 << 2'h2;
  assign T29 = io_in_1 & 2'h3;
  assign T30 = T49 & T31;
  assign T31 = ~ T32;
  assign T32 = 5'hc;
  assign T49 = {2'h0, T33};
  assign T33 = T36 | T50;
  assign T50 = {1'h0, T34};
  assign T34 = T35 << 1'h0;
  assign T35 = io_in_0 & 2'h3;
  assign T36 = 3'h0 & T37;
  assign T37 = ~ T38;
  assign T38 = 3'h3;
  assign io_out = VwireFlatBlackBox_out;
  vwire #(.W(2),.L(3)) VwireFlatBlackBox(
       .in( T45 ),
       .en( T39 ),
       .out( VwireFlatBlackBox_out )
  );
endmodule

module Vwire3BB(
    input [1:0] io_in_2,
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    input  io_en_2,
    input  io_en_1,
    input  io_en_0,
    output[1:0] io_out
);

  wire[1:0] VwireBlackBox_io_out;


  assign io_out = VwireBlackBox_io_out;
  VwireBlackBox_1 VwireBlackBox(
       .io_in_2( io_in_2 ),
       .io_in_1( io_in_1 ),
       .io_in_0( io_in_0 ),
       .io_en_2( io_en_2 ),
       .io_en_1( io_en_1 ),
       .io_en_0( io_en_0 ),
       .io_out( VwireBlackBox_io_out )
  );
endmodule

module Vwire_1(
    input [1:0] io_in_2,
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    input  io_en_2,
    input  io_en_1,
    input  io_en_0,
    output[1:0] io_out
);

  wire[1:0] Vwire3BB_io_out;


  assign io_out = Vwire3BB_io_out;
  Vwire3BB Vwire3BB(
       .io_in_2( io_in_2 ),
       .io_in_1( io_in_1 ),
       .io_in_0( io_in_0 ),
       .io_en_2( io_en_2 ),
       .io_en_1( io_en_1 ),
       .io_en_0( io_en_0 ),
       .io_out( Vwire3BB_io_out )
  );
endmodule

module VwireBlackBox_2(
    input [1:0] io_in_3,
    input [1:0] io_in_2,
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    input  io_en_3,
    input  io_en_2,
    input  io_en_1,
    input  io_en_0,
    output[1:0] io_out
);

  wire[3:0] T52;
  wire[4:0] T0;
  wire[4:0] T1;
  wire[4:0] T2;
  wire[4:0] T53;
  wire T3;
  wire T4;
  wire[4:0] T5;
  wire[4:0] T6;
  wire[4:0] T54;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T55;
  wire T10;
  wire T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T56;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T57;
  wire T17;
  wire T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T58;
  wire[1:0] T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire[1:0] T59;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire[7:0] T60;
  wire[8:0] T28;
  wire[8:0] T61;
  wire[7:0] T29;
  wire[1:0] T30;
  wire[8:0] T31;
  wire[8:0] T32;
  wire[8:0] T33;
  wire[8:0] T62;
  wire[6:0] T34;
  wire[6:0] T63;
  wire[5:0] T35;
  wire[1:0] T36;
  wire[6:0] T37;
  wire[6:0] T38;
  wire[6:0] T39;
  wire[6:0] T64;
  wire[4:0] T40;
  wire[4:0] T65;
  wire[3:0] T41;
  wire[1:0] T42;
  wire[4:0] T43;
  wire[4:0] T44;
  wire[4:0] T45;
  wire[4:0] T66;
  wire[2:0] T46;
  wire[2:0] T67;
  wire[1:0] T47;
  wire[1:0] T48;
  wire[2:0] T49;
  wire[2:0] T50;
  wire[2:0] T51;
  wire[1:0] VwireFlatBlackBox_out;


  assign T52 = T0[2'h3:1'h0];
  assign T0 = T5 | T1;
  assign T1 = T53 & T2;
  assign T2 = 5'h8;
  assign T53 = T3 ? 5'h1f : 5'h0;
  assign T3 = T4;
  assign T4 = io_en_3;
  assign T5 = T54 & T6;
  assign T6 = ~ T2;
  assign T54 = {1'h0, T7};
  assign T7 = T12 | T8;
  assign T8 = T55 & T9;
  assign T9 = 4'h4;
  assign T55 = T10 ? 4'hf : 4'h0;
  assign T10 = T11;
  assign T11 = io_en_2;
  assign T12 = T56 & T13;
  assign T13 = ~ T9;
  assign T56 = {1'h0, T14};
  assign T14 = T19 | T15;
  assign T15 = T57 & T16;
  assign T16 = 3'h2;
  assign T57 = T17 ? 3'h7 : 3'h0;
  assign T17 = T18;
  assign T18 = io_en_1;
  assign T19 = T58 & T20;
  assign T20 = ~ T16;
  assign T58 = {1'h0, T21};
  assign T21 = T26 | T22;
  assign T22 = T59 & T23;
  assign T23 = 2'h1;
  assign T59 = T24 ? 2'h3 : 2'h0;
  assign T24 = T25;
  assign T25 = io_en_0;
  assign T26 = 2'h0 & T27;
  assign T27 = ~ T23;
  assign T60 = T28[3'h7:1'h0];
  assign T28 = T31 | T61;
  assign T61 = {1'h0, T29};
  assign T29 = T30 << 3'h6;
  assign T30 = io_in_3 & 2'h3;
  assign T31 = T62 & T32;
  assign T32 = ~ T33;
  assign T33 = 9'hc0;
  assign T62 = {2'h0, T34};
  assign T34 = T37 | T63;
  assign T63 = {1'h0, T35};
  assign T35 = T36 << 3'h4;
  assign T36 = io_in_2 & 2'h3;
  assign T37 = T64 & T38;
  assign T38 = ~ T39;
  assign T39 = 7'h30;
  assign T64 = {2'h0, T40};
  assign T40 = T43 | T65;
  assign T65 = {1'h0, T41};
  assign T41 = T42 << 2'h2;
  assign T42 = io_in_1 & 2'h3;
  assign T43 = T66 & T44;
  assign T44 = ~ T45;
  assign T45 = 5'hc;
  assign T66 = {2'h0, T46};
  assign T46 = T49 | T67;
  assign T67 = {1'h0, T47};
  assign T47 = T48 << 1'h0;
  assign T48 = io_in_0 & 2'h3;
  assign T49 = 3'h0 & T50;
  assign T50 = ~ T51;
  assign T51 = 3'h3;
  assign io_out = VwireFlatBlackBox_out;
  vwire #(.W(2),.L(4)) VwireFlatBlackBox(
       .in( T60 ),
       .en( T52 ),
       .out( VwireFlatBlackBox_out )
  );
endmodule

module Vwire4BB(
    input [1:0] io_in_3,
    input [1:0] io_in_2,
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    input  io_en_3,
    input  io_en_2,
    input  io_en_1,
    input  io_en_0,
    output[1:0] io_out
);

  wire[1:0] VwireBlackBox_io_out;


  assign io_out = VwireBlackBox_io_out;
  VwireBlackBox_2 VwireBlackBox(
       .io_in_3( io_in_3 ),
       .io_in_2( io_in_2 ),
       .io_in_1( io_in_1 ),
       .io_in_0( io_in_0 ),
       .io_en_3( io_en_3 ),
       .io_en_2( io_en_2 ),
       .io_en_1( io_en_1 ),
       .io_en_0( io_en_0 ),
       .io_out( VwireBlackBox_io_out )
  );
endmodule

module Vwire_2(
    input [1:0] io_in_3,
    input [1:0] io_in_2,
    input [1:0] io_in_1,
    input [1:0] io_in_0,
    input  io_en_3,
    input  io_en_2,
    input  io_en_1,
    input  io_en_0,
    output[1:0] io_out
);

  wire[1:0] Vwire4BB_io_out;


  assign io_out = Vwire4BB_io_out;
  Vwire4BB Vwire4BB(
       .io_in_3( io_in_3 ),
       .io_in_2( io_in_2 ),
       .io_in_1( io_in_1 ),
       .io_in_0( io_in_0 ),
       .io_en_3( io_en_3 ),
       .io_en_2( io_en_2 ),
       .io_en_1( io_en_1 ),
       .io_en_0( io_en_0 ),
       .io_out( Vwire4BB_io_out )
  );
endmodule

module VwireModule(
    input [1:0] io_VwirePorts_3_22_15_in,
    input  io_VwirePorts_3_22_15_en,
    output[1:0] io_VwirePorts_3_22_15_out,
    input [1:0] io_VwirePorts_3_22_14_in,
    input  io_VwirePorts_3_22_14_en,
    output[1:0] io_VwirePorts_3_22_14_out,
    input [1:0] io_VwirePorts_3_22_13_in,
    input  io_VwirePorts_3_22_13_en,
    output[1:0] io_VwirePorts_3_22_13_out,
    input [1:0] io_VwirePorts_3_22_12_in,
    input  io_VwirePorts_3_22_12_en,
    output[1:0] io_VwirePorts_3_22_12_out,
    input [1:0] io_VwirePorts_3_22_11_in,
    input  io_VwirePorts_3_22_11_en,
    output[1:0] io_VwirePorts_3_22_11_out,
    input [1:0] io_VwirePorts_3_22_10_in,
    input  io_VwirePorts_3_22_10_en,
    output[1:0] io_VwirePorts_3_22_10_out,
    input [1:0] io_VwirePorts_3_22_9_in,
    input  io_VwirePorts_3_22_9_en,
    output[1:0] io_VwirePorts_3_22_9_out,
    input [1:0] io_VwirePorts_3_22_8_in,
    input  io_VwirePorts_3_22_8_en,
    output[1:0] io_VwirePorts_3_22_8_out,
    input [1:0] io_VwirePorts_3_22_7_in,
    input  io_VwirePorts_3_22_7_en,
    output[1:0] io_VwirePorts_3_22_7_out,
    input [1:0] io_VwirePorts_3_22_6_in,
    input  io_VwirePorts_3_22_6_en,
    output[1:0] io_VwirePorts_3_22_6_out,
    input [1:0] io_VwirePorts_3_22_5_in,
    input  io_VwirePorts_3_22_5_en,
    output[1:0] io_VwirePorts_3_22_5_out,
    input [1:0] io_VwirePorts_3_22_4_in,
    input  io_VwirePorts_3_22_4_en,
    output[1:0] io_VwirePorts_3_22_4_out,
    input [1:0] io_VwirePorts_3_22_3_in,
    input  io_VwirePorts_3_22_3_en,
    output[1:0] io_VwirePorts_3_22_3_out,
    input [1:0] io_VwirePorts_3_22_2_in,
    input  io_VwirePorts_3_22_2_en,
    output[1:0] io_VwirePorts_3_22_2_out,
    input [1:0] io_VwirePorts_3_22_1_in,
    input  io_VwirePorts_3_22_1_en,
    output[1:0] io_VwirePorts_3_22_1_out,
    input [1:0] io_VwirePorts_3_22_0_in,
    input  io_VwirePorts_3_22_0_en,
    output[1:0] io_VwirePorts_3_22_0_out,
    input [1:0] io_VwirePorts_3_21_15_in,
    input  io_VwirePorts_3_21_15_en,
    output[1:0] io_VwirePorts_3_21_15_out,
    input [1:0] io_VwirePorts_3_21_14_in,
    input  io_VwirePorts_3_21_14_en,
    output[1:0] io_VwirePorts_3_21_14_out,
    input [1:0] io_VwirePorts_3_21_13_in,
    input  io_VwirePorts_3_21_13_en,
    output[1:0] io_VwirePorts_3_21_13_out,
    input [1:0] io_VwirePorts_3_21_12_in,
    input  io_VwirePorts_3_21_12_en,
    output[1:0] io_VwirePorts_3_21_12_out,
    input [1:0] io_VwirePorts_3_21_11_in,
    input  io_VwirePorts_3_21_11_en,
    output[1:0] io_VwirePorts_3_21_11_out,
    input [1:0] io_VwirePorts_3_21_10_in,
    input  io_VwirePorts_3_21_10_en,
    output[1:0] io_VwirePorts_3_21_10_out,
    input [1:0] io_VwirePorts_3_21_9_in,
    input  io_VwirePorts_3_21_9_en,
    output[1:0] io_VwirePorts_3_21_9_out,
    input [1:0] io_VwirePorts_3_21_8_in,
    input  io_VwirePorts_3_21_8_en,
    output[1:0] io_VwirePorts_3_21_8_out,
    input [1:0] io_VwirePorts_3_21_7_in,
    input  io_VwirePorts_3_21_7_en,
    output[1:0] io_VwirePorts_3_21_7_out,
    input [1:0] io_VwirePorts_3_21_6_in,
    input  io_VwirePorts_3_21_6_en,
    output[1:0] io_VwirePorts_3_21_6_out,
    input [1:0] io_VwirePorts_3_21_5_in,
    input  io_VwirePorts_3_21_5_en,
    output[1:0] io_VwirePorts_3_21_5_out,
    input [1:0] io_VwirePorts_3_21_4_in,
    input  io_VwirePorts_3_21_4_en,
    output[1:0] io_VwirePorts_3_21_4_out,
    input [1:0] io_VwirePorts_3_21_3_in,
    input  io_VwirePorts_3_21_3_en,
    output[1:0] io_VwirePorts_3_21_3_out,
    input [1:0] io_VwirePorts_3_21_2_in,
    input  io_VwirePorts_3_21_2_en,
    output[1:0] io_VwirePorts_3_21_2_out,
    input [1:0] io_VwirePorts_3_21_1_in,
    input  io_VwirePorts_3_21_1_en,
    output[1:0] io_VwirePorts_3_21_1_out,
    input [1:0] io_VwirePorts_3_21_0_in,
    input  io_VwirePorts_3_21_0_en,
    output[1:0] io_VwirePorts_3_21_0_out,
    input [1:0] io_VwirePorts_3_20_15_in,
    input  io_VwirePorts_3_20_15_en,
    output[1:0] io_VwirePorts_3_20_15_out,
    input [1:0] io_VwirePorts_3_20_14_in,
    input  io_VwirePorts_3_20_14_en,
    output[1:0] io_VwirePorts_3_20_14_out,
    input [1:0] io_VwirePorts_3_20_13_in,
    input  io_VwirePorts_3_20_13_en,
    output[1:0] io_VwirePorts_3_20_13_out,
    input [1:0] io_VwirePorts_3_20_12_in,
    input  io_VwirePorts_3_20_12_en,
    output[1:0] io_VwirePorts_3_20_12_out,
    input [1:0] io_VwirePorts_3_20_11_in,
    input  io_VwirePorts_3_20_11_en,
    output[1:0] io_VwirePorts_3_20_11_out,
    input [1:0] io_VwirePorts_3_20_10_in,
    input  io_VwirePorts_3_20_10_en,
    output[1:0] io_VwirePorts_3_20_10_out,
    input [1:0] io_VwirePorts_3_20_9_in,
    input  io_VwirePorts_3_20_9_en,
    output[1:0] io_VwirePorts_3_20_9_out,
    input [1:0] io_VwirePorts_3_20_8_in,
    input  io_VwirePorts_3_20_8_en,
    output[1:0] io_VwirePorts_3_20_8_out,
    input [1:0] io_VwirePorts_3_20_7_in,
    input  io_VwirePorts_3_20_7_en,
    output[1:0] io_VwirePorts_3_20_7_out,
    input [1:0] io_VwirePorts_3_20_6_in,
    input  io_VwirePorts_3_20_6_en,
    output[1:0] io_VwirePorts_3_20_6_out,
    input [1:0] io_VwirePorts_3_20_5_in,
    input  io_VwirePorts_3_20_5_en,
    output[1:0] io_VwirePorts_3_20_5_out,
    input [1:0] io_VwirePorts_3_20_4_in,
    input  io_VwirePorts_3_20_4_en,
    output[1:0] io_VwirePorts_3_20_4_out,
    input [1:0] io_VwirePorts_3_20_3_in,
    input  io_VwirePorts_3_20_3_en,
    output[1:0] io_VwirePorts_3_20_3_out,
    input [1:0] io_VwirePorts_3_20_2_in,
    input  io_VwirePorts_3_20_2_en,
    output[1:0] io_VwirePorts_3_20_2_out,
    input [1:0] io_VwirePorts_3_20_1_in,
    input  io_VwirePorts_3_20_1_en,
    output[1:0] io_VwirePorts_3_20_1_out,
    input [1:0] io_VwirePorts_3_20_0_in,
    input  io_VwirePorts_3_20_0_en,
    output[1:0] io_VwirePorts_3_20_0_out,
    input [1:0] io_VwirePorts_3_19_15_in,
    input  io_VwirePorts_3_19_15_en,
    output[1:0] io_VwirePorts_3_19_15_out,
    input [1:0] io_VwirePorts_3_19_14_in,
    input  io_VwirePorts_3_19_14_en,
    output[1:0] io_VwirePorts_3_19_14_out,
    input [1:0] io_VwirePorts_3_19_13_in,
    input  io_VwirePorts_3_19_13_en,
    output[1:0] io_VwirePorts_3_19_13_out,
    input [1:0] io_VwirePorts_3_19_12_in,
    input  io_VwirePorts_3_19_12_en,
    output[1:0] io_VwirePorts_3_19_12_out,
    input [1:0] io_VwirePorts_3_19_11_in,
    input  io_VwirePorts_3_19_11_en,
    output[1:0] io_VwirePorts_3_19_11_out,
    input [1:0] io_VwirePorts_3_19_10_in,
    input  io_VwirePorts_3_19_10_en,
    output[1:0] io_VwirePorts_3_19_10_out,
    input [1:0] io_VwirePorts_3_19_9_in,
    input  io_VwirePorts_3_19_9_en,
    output[1:0] io_VwirePorts_3_19_9_out,
    input [1:0] io_VwirePorts_3_19_8_in,
    input  io_VwirePorts_3_19_8_en,
    output[1:0] io_VwirePorts_3_19_8_out,
    input [1:0] io_VwirePorts_3_19_7_in,
    input  io_VwirePorts_3_19_7_en,
    output[1:0] io_VwirePorts_3_19_7_out,
    input [1:0] io_VwirePorts_3_19_6_in,
    input  io_VwirePorts_3_19_6_en,
    output[1:0] io_VwirePorts_3_19_6_out,
    input [1:0] io_VwirePorts_3_19_5_in,
    input  io_VwirePorts_3_19_5_en,
    output[1:0] io_VwirePorts_3_19_5_out,
    input [1:0] io_VwirePorts_3_19_4_in,
    input  io_VwirePorts_3_19_4_en,
    output[1:0] io_VwirePorts_3_19_4_out,
    input [1:0] io_VwirePorts_3_19_3_in,
    input  io_VwirePorts_3_19_3_en,
    output[1:0] io_VwirePorts_3_19_3_out,
    input [1:0] io_VwirePorts_3_19_2_in,
    input  io_VwirePorts_3_19_2_en,
    output[1:0] io_VwirePorts_3_19_2_out,
    input [1:0] io_VwirePorts_3_19_1_in,
    input  io_VwirePorts_3_19_1_en,
    output[1:0] io_VwirePorts_3_19_1_out,
    input [1:0] io_VwirePorts_3_19_0_in,
    input  io_VwirePorts_3_19_0_en,
    output[1:0] io_VwirePorts_3_19_0_out,
    input [1:0] io_VwirePorts_3_18_15_in,
    input  io_VwirePorts_3_18_15_en,
    output[1:0] io_VwirePorts_3_18_15_out,
    input [1:0] io_VwirePorts_3_18_14_in,
    input  io_VwirePorts_3_18_14_en,
    output[1:0] io_VwirePorts_3_18_14_out,
    input [1:0] io_VwirePorts_3_18_13_in,
    input  io_VwirePorts_3_18_13_en,
    output[1:0] io_VwirePorts_3_18_13_out,
    input [1:0] io_VwirePorts_3_18_12_in,
    input  io_VwirePorts_3_18_12_en,
    output[1:0] io_VwirePorts_3_18_12_out,
    input [1:0] io_VwirePorts_3_18_11_in,
    input  io_VwirePorts_3_18_11_en,
    output[1:0] io_VwirePorts_3_18_11_out,
    input [1:0] io_VwirePorts_3_18_10_in,
    input  io_VwirePorts_3_18_10_en,
    output[1:0] io_VwirePorts_3_18_10_out,
    input [1:0] io_VwirePorts_3_18_9_in,
    input  io_VwirePorts_3_18_9_en,
    output[1:0] io_VwirePorts_3_18_9_out,
    input [1:0] io_VwirePorts_3_18_8_in,
    input  io_VwirePorts_3_18_8_en,
    output[1:0] io_VwirePorts_3_18_8_out,
    input [1:0] io_VwirePorts_3_18_7_in,
    input  io_VwirePorts_3_18_7_en,
    output[1:0] io_VwirePorts_3_18_7_out,
    input [1:0] io_VwirePorts_3_18_6_in,
    input  io_VwirePorts_3_18_6_en,
    output[1:0] io_VwirePorts_3_18_6_out,
    input [1:0] io_VwirePorts_3_18_5_in,
    input  io_VwirePorts_3_18_5_en,
    output[1:0] io_VwirePorts_3_18_5_out,
    input [1:0] io_VwirePorts_3_18_4_in,
    input  io_VwirePorts_3_18_4_en,
    output[1:0] io_VwirePorts_3_18_4_out,
    input [1:0] io_VwirePorts_3_18_3_in,
    input  io_VwirePorts_3_18_3_en,
    output[1:0] io_VwirePorts_3_18_3_out,
    input [1:0] io_VwirePorts_3_18_2_in,
    input  io_VwirePorts_3_18_2_en,
    output[1:0] io_VwirePorts_3_18_2_out,
    input [1:0] io_VwirePorts_3_18_1_in,
    input  io_VwirePorts_3_18_1_en,
    output[1:0] io_VwirePorts_3_18_1_out,
    input [1:0] io_VwirePorts_3_18_0_in,
    input  io_VwirePorts_3_18_0_en,
    output[1:0] io_VwirePorts_3_18_0_out,
    input [1:0] io_VwirePorts_3_17_15_in,
    input  io_VwirePorts_3_17_15_en,
    output[1:0] io_VwirePorts_3_17_15_out,
    input [1:0] io_VwirePorts_3_17_14_in,
    input  io_VwirePorts_3_17_14_en,
    output[1:0] io_VwirePorts_3_17_14_out,
    input [1:0] io_VwirePorts_3_17_13_in,
    input  io_VwirePorts_3_17_13_en,
    output[1:0] io_VwirePorts_3_17_13_out,
    input [1:0] io_VwirePorts_3_17_12_in,
    input  io_VwirePorts_3_17_12_en,
    output[1:0] io_VwirePorts_3_17_12_out,
    input [1:0] io_VwirePorts_3_17_11_in,
    input  io_VwirePorts_3_17_11_en,
    output[1:0] io_VwirePorts_3_17_11_out,
    input [1:0] io_VwirePorts_3_17_10_in,
    input  io_VwirePorts_3_17_10_en,
    output[1:0] io_VwirePorts_3_17_10_out,
    input [1:0] io_VwirePorts_3_17_9_in,
    input  io_VwirePorts_3_17_9_en,
    output[1:0] io_VwirePorts_3_17_9_out,
    input [1:0] io_VwirePorts_3_17_8_in,
    input  io_VwirePorts_3_17_8_en,
    output[1:0] io_VwirePorts_3_17_8_out,
    input [1:0] io_VwirePorts_3_17_7_in,
    input  io_VwirePorts_3_17_7_en,
    output[1:0] io_VwirePorts_3_17_7_out,
    input [1:0] io_VwirePorts_3_17_6_in,
    input  io_VwirePorts_3_17_6_en,
    output[1:0] io_VwirePorts_3_17_6_out,
    input [1:0] io_VwirePorts_3_17_5_in,
    input  io_VwirePorts_3_17_5_en,
    output[1:0] io_VwirePorts_3_17_5_out,
    input [1:0] io_VwirePorts_3_17_4_in,
    input  io_VwirePorts_3_17_4_en,
    output[1:0] io_VwirePorts_3_17_4_out,
    input [1:0] io_VwirePorts_3_17_3_in,
    input  io_VwirePorts_3_17_3_en,
    output[1:0] io_VwirePorts_3_17_3_out,
    input [1:0] io_VwirePorts_3_17_2_in,
    input  io_VwirePorts_3_17_2_en,
    output[1:0] io_VwirePorts_3_17_2_out,
    input [1:0] io_VwirePorts_3_17_1_in,
    input  io_VwirePorts_3_17_1_en,
    output[1:0] io_VwirePorts_3_17_1_out,
    input [1:0] io_VwirePorts_3_17_0_in,
    input  io_VwirePorts_3_17_0_en,
    output[1:0] io_VwirePorts_3_17_0_out,
    input [1:0] io_VwirePorts_3_16_15_in,
    input  io_VwirePorts_3_16_15_en,
    output[1:0] io_VwirePorts_3_16_15_out,
    input [1:0] io_VwirePorts_3_16_14_in,
    input  io_VwirePorts_3_16_14_en,
    output[1:0] io_VwirePorts_3_16_14_out,
    input [1:0] io_VwirePorts_3_16_13_in,
    input  io_VwirePorts_3_16_13_en,
    output[1:0] io_VwirePorts_3_16_13_out,
    input [1:0] io_VwirePorts_3_16_12_in,
    input  io_VwirePorts_3_16_12_en,
    output[1:0] io_VwirePorts_3_16_12_out,
    input [1:0] io_VwirePorts_3_16_11_in,
    input  io_VwirePorts_3_16_11_en,
    output[1:0] io_VwirePorts_3_16_11_out,
    input [1:0] io_VwirePorts_3_16_10_in,
    input  io_VwirePorts_3_16_10_en,
    output[1:0] io_VwirePorts_3_16_10_out,
    input [1:0] io_VwirePorts_3_16_9_in,
    input  io_VwirePorts_3_16_9_en,
    output[1:0] io_VwirePorts_3_16_9_out,
    input [1:0] io_VwirePorts_3_16_8_in,
    input  io_VwirePorts_3_16_8_en,
    output[1:0] io_VwirePorts_3_16_8_out,
    input [1:0] io_VwirePorts_3_16_7_in,
    input  io_VwirePorts_3_16_7_en,
    output[1:0] io_VwirePorts_3_16_7_out,
    input [1:0] io_VwirePorts_3_16_6_in,
    input  io_VwirePorts_3_16_6_en,
    output[1:0] io_VwirePorts_3_16_6_out,
    input [1:0] io_VwirePorts_3_16_5_in,
    input  io_VwirePorts_3_16_5_en,
    output[1:0] io_VwirePorts_3_16_5_out,
    input [1:0] io_VwirePorts_3_16_4_in,
    input  io_VwirePorts_3_16_4_en,
    output[1:0] io_VwirePorts_3_16_4_out,
    input [1:0] io_VwirePorts_3_16_3_in,
    input  io_VwirePorts_3_16_3_en,
    output[1:0] io_VwirePorts_3_16_3_out,
    input [1:0] io_VwirePorts_3_16_2_in,
    input  io_VwirePorts_3_16_2_en,
    output[1:0] io_VwirePorts_3_16_2_out,
    input [1:0] io_VwirePorts_3_16_1_in,
    input  io_VwirePorts_3_16_1_en,
    output[1:0] io_VwirePorts_3_16_1_out,
    input [1:0] io_VwirePorts_3_16_0_in,
    input  io_VwirePorts_3_16_0_en,
    output[1:0] io_VwirePorts_3_16_0_out,
    input [1:0] io_VwirePorts_3_15_15_in,
    input  io_VwirePorts_3_15_15_en,
    output[1:0] io_VwirePorts_3_15_15_out,
    input [1:0] io_VwirePorts_3_15_14_in,
    input  io_VwirePorts_3_15_14_en,
    output[1:0] io_VwirePorts_3_15_14_out,
    input [1:0] io_VwirePorts_3_15_13_in,
    input  io_VwirePorts_3_15_13_en,
    output[1:0] io_VwirePorts_3_15_13_out,
    input [1:0] io_VwirePorts_3_15_12_in,
    input  io_VwirePorts_3_15_12_en,
    output[1:0] io_VwirePorts_3_15_12_out,
    input [1:0] io_VwirePorts_3_15_11_in,
    input  io_VwirePorts_3_15_11_en,
    output[1:0] io_VwirePorts_3_15_11_out,
    input [1:0] io_VwirePorts_3_15_10_in,
    input  io_VwirePorts_3_15_10_en,
    output[1:0] io_VwirePorts_3_15_10_out,
    input [1:0] io_VwirePorts_3_15_9_in,
    input  io_VwirePorts_3_15_9_en,
    output[1:0] io_VwirePorts_3_15_9_out,
    input [1:0] io_VwirePorts_3_15_8_in,
    input  io_VwirePorts_3_15_8_en,
    output[1:0] io_VwirePorts_3_15_8_out,
    input [1:0] io_VwirePorts_3_15_7_in,
    input  io_VwirePorts_3_15_7_en,
    output[1:0] io_VwirePorts_3_15_7_out,
    input [1:0] io_VwirePorts_3_15_6_in,
    input  io_VwirePorts_3_15_6_en,
    output[1:0] io_VwirePorts_3_15_6_out,
    input [1:0] io_VwirePorts_3_15_5_in,
    input  io_VwirePorts_3_15_5_en,
    output[1:0] io_VwirePorts_3_15_5_out,
    input [1:0] io_VwirePorts_3_15_4_in,
    input  io_VwirePorts_3_15_4_en,
    output[1:0] io_VwirePorts_3_15_4_out,
    input [1:0] io_VwirePorts_3_15_3_in,
    input  io_VwirePorts_3_15_3_en,
    output[1:0] io_VwirePorts_3_15_3_out,
    input [1:0] io_VwirePorts_3_15_2_in,
    input  io_VwirePorts_3_15_2_en,
    output[1:0] io_VwirePorts_3_15_2_out,
    input [1:0] io_VwirePorts_3_15_1_in,
    input  io_VwirePorts_3_15_1_en,
    output[1:0] io_VwirePorts_3_15_1_out,
    input [1:0] io_VwirePorts_3_15_0_in,
    input  io_VwirePorts_3_15_0_en,
    output[1:0] io_VwirePorts_3_15_0_out,
    input [1:0] io_VwirePorts_3_14_15_in,
    input  io_VwirePorts_3_14_15_en,
    output[1:0] io_VwirePorts_3_14_15_out,
    input [1:0] io_VwirePorts_3_14_14_in,
    input  io_VwirePorts_3_14_14_en,
    output[1:0] io_VwirePorts_3_14_14_out,
    input [1:0] io_VwirePorts_3_14_13_in,
    input  io_VwirePorts_3_14_13_en,
    output[1:0] io_VwirePorts_3_14_13_out,
    input [1:0] io_VwirePorts_3_14_12_in,
    input  io_VwirePorts_3_14_12_en,
    output[1:0] io_VwirePorts_3_14_12_out,
    input [1:0] io_VwirePorts_3_14_11_in,
    input  io_VwirePorts_3_14_11_en,
    output[1:0] io_VwirePorts_3_14_11_out,
    input [1:0] io_VwirePorts_3_14_10_in,
    input  io_VwirePorts_3_14_10_en,
    output[1:0] io_VwirePorts_3_14_10_out,
    input [1:0] io_VwirePorts_3_14_9_in,
    input  io_VwirePorts_3_14_9_en,
    output[1:0] io_VwirePorts_3_14_9_out,
    input [1:0] io_VwirePorts_3_14_8_in,
    input  io_VwirePorts_3_14_8_en,
    output[1:0] io_VwirePorts_3_14_8_out,
    input [1:0] io_VwirePorts_3_14_7_in,
    input  io_VwirePorts_3_14_7_en,
    output[1:0] io_VwirePorts_3_14_7_out,
    input [1:0] io_VwirePorts_3_14_6_in,
    input  io_VwirePorts_3_14_6_en,
    output[1:0] io_VwirePorts_3_14_6_out,
    input [1:0] io_VwirePorts_3_14_5_in,
    input  io_VwirePorts_3_14_5_en,
    output[1:0] io_VwirePorts_3_14_5_out,
    input [1:0] io_VwirePorts_3_14_4_in,
    input  io_VwirePorts_3_14_4_en,
    output[1:0] io_VwirePorts_3_14_4_out,
    input [1:0] io_VwirePorts_3_14_3_in,
    input  io_VwirePorts_3_14_3_en,
    output[1:0] io_VwirePorts_3_14_3_out,
    input [1:0] io_VwirePorts_3_14_2_in,
    input  io_VwirePorts_3_14_2_en,
    output[1:0] io_VwirePorts_3_14_2_out,
    input [1:0] io_VwirePorts_3_14_1_in,
    input  io_VwirePorts_3_14_1_en,
    output[1:0] io_VwirePorts_3_14_1_out,
    input [1:0] io_VwirePorts_3_14_0_in,
    input  io_VwirePorts_3_14_0_en,
    output[1:0] io_VwirePorts_3_14_0_out,
    input [1:0] io_VwirePorts_3_13_15_in,
    input  io_VwirePorts_3_13_15_en,
    output[1:0] io_VwirePorts_3_13_15_out,
    input [1:0] io_VwirePorts_3_13_14_in,
    input  io_VwirePorts_3_13_14_en,
    output[1:0] io_VwirePorts_3_13_14_out,
    input [1:0] io_VwirePorts_3_13_13_in,
    input  io_VwirePorts_3_13_13_en,
    output[1:0] io_VwirePorts_3_13_13_out,
    input [1:0] io_VwirePorts_3_13_12_in,
    input  io_VwirePorts_3_13_12_en,
    output[1:0] io_VwirePorts_3_13_12_out,
    input [1:0] io_VwirePorts_3_13_11_in,
    input  io_VwirePorts_3_13_11_en,
    output[1:0] io_VwirePorts_3_13_11_out,
    input [1:0] io_VwirePorts_3_13_10_in,
    input  io_VwirePorts_3_13_10_en,
    output[1:0] io_VwirePorts_3_13_10_out,
    input [1:0] io_VwirePorts_3_13_9_in,
    input  io_VwirePorts_3_13_9_en,
    output[1:0] io_VwirePorts_3_13_9_out,
    input [1:0] io_VwirePorts_3_13_8_in,
    input  io_VwirePorts_3_13_8_en,
    output[1:0] io_VwirePorts_3_13_8_out,
    input [1:0] io_VwirePorts_3_13_7_in,
    input  io_VwirePorts_3_13_7_en,
    output[1:0] io_VwirePorts_3_13_7_out,
    input [1:0] io_VwirePorts_3_13_6_in,
    input  io_VwirePorts_3_13_6_en,
    output[1:0] io_VwirePorts_3_13_6_out,
    input [1:0] io_VwirePorts_3_13_5_in,
    input  io_VwirePorts_3_13_5_en,
    output[1:0] io_VwirePorts_3_13_5_out,
    input [1:0] io_VwirePorts_3_13_4_in,
    input  io_VwirePorts_3_13_4_en,
    output[1:0] io_VwirePorts_3_13_4_out,
    input [1:0] io_VwirePorts_3_13_3_in,
    input  io_VwirePorts_3_13_3_en,
    output[1:0] io_VwirePorts_3_13_3_out,
    input [1:0] io_VwirePorts_3_13_2_in,
    input  io_VwirePorts_3_13_2_en,
    output[1:0] io_VwirePorts_3_13_2_out,
    input [1:0] io_VwirePorts_3_13_1_in,
    input  io_VwirePorts_3_13_1_en,
    output[1:0] io_VwirePorts_3_13_1_out,
    input [1:0] io_VwirePorts_3_13_0_in,
    input  io_VwirePorts_3_13_0_en,
    output[1:0] io_VwirePorts_3_13_0_out,
    input [1:0] io_VwirePorts_3_12_15_in,
    input  io_VwirePorts_3_12_15_en,
    output[1:0] io_VwirePorts_3_12_15_out,
    input [1:0] io_VwirePorts_3_12_14_in,
    input  io_VwirePorts_3_12_14_en,
    output[1:0] io_VwirePorts_3_12_14_out,
    input [1:0] io_VwirePorts_3_12_13_in,
    input  io_VwirePorts_3_12_13_en,
    output[1:0] io_VwirePorts_3_12_13_out,
    input [1:0] io_VwirePorts_3_12_12_in,
    input  io_VwirePorts_3_12_12_en,
    output[1:0] io_VwirePorts_3_12_12_out,
    input [1:0] io_VwirePorts_3_12_11_in,
    input  io_VwirePorts_3_12_11_en,
    output[1:0] io_VwirePorts_3_12_11_out,
    input [1:0] io_VwirePorts_3_12_10_in,
    input  io_VwirePorts_3_12_10_en,
    output[1:0] io_VwirePorts_3_12_10_out,
    input [1:0] io_VwirePorts_3_12_9_in,
    input  io_VwirePorts_3_12_9_en,
    output[1:0] io_VwirePorts_3_12_9_out,
    input [1:0] io_VwirePorts_3_12_8_in,
    input  io_VwirePorts_3_12_8_en,
    output[1:0] io_VwirePorts_3_12_8_out,
    input [1:0] io_VwirePorts_3_12_7_in,
    input  io_VwirePorts_3_12_7_en,
    output[1:0] io_VwirePorts_3_12_7_out,
    input [1:0] io_VwirePorts_3_12_6_in,
    input  io_VwirePorts_3_12_6_en,
    output[1:0] io_VwirePorts_3_12_6_out,
    input [1:0] io_VwirePorts_3_12_5_in,
    input  io_VwirePorts_3_12_5_en,
    output[1:0] io_VwirePorts_3_12_5_out,
    input [1:0] io_VwirePorts_3_12_4_in,
    input  io_VwirePorts_3_12_4_en,
    output[1:0] io_VwirePorts_3_12_4_out,
    input [1:0] io_VwirePorts_3_12_3_in,
    input  io_VwirePorts_3_12_3_en,
    output[1:0] io_VwirePorts_3_12_3_out,
    input [1:0] io_VwirePorts_3_12_2_in,
    input  io_VwirePorts_3_12_2_en,
    output[1:0] io_VwirePorts_3_12_2_out,
    input [1:0] io_VwirePorts_3_12_1_in,
    input  io_VwirePorts_3_12_1_en,
    output[1:0] io_VwirePorts_3_12_1_out,
    input [1:0] io_VwirePorts_3_12_0_in,
    input  io_VwirePorts_3_12_0_en,
    output[1:0] io_VwirePorts_3_12_0_out,
    input [1:0] io_VwirePorts_3_11_15_in,
    input  io_VwirePorts_3_11_15_en,
    output[1:0] io_VwirePorts_3_11_15_out,
    input [1:0] io_VwirePorts_3_11_14_in,
    input  io_VwirePorts_3_11_14_en,
    output[1:0] io_VwirePorts_3_11_14_out,
    input [1:0] io_VwirePorts_3_11_13_in,
    input  io_VwirePorts_3_11_13_en,
    output[1:0] io_VwirePorts_3_11_13_out,
    input [1:0] io_VwirePorts_3_11_12_in,
    input  io_VwirePorts_3_11_12_en,
    output[1:0] io_VwirePorts_3_11_12_out,
    input [1:0] io_VwirePorts_3_11_11_in,
    input  io_VwirePorts_3_11_11_en,
    output[1:0] io_VwirePorts_3_11_11_out,
    input [1:0] io_VwirePorts_3_11_10_in,
    input  io_VwirePorts_3_11_10_en,
    output[1:0] io_VwirePorts_3_11_10_out,
    input [1:0] io_VwirePorts_3_11_9_in,
    input  io_VwirePorts_3_11_9_en,
    output[1:0] io_VwirePorts_3_11_9_out,
    input [1:0] io_VwirePorts_3_11_8_in,
    input  io_VwirePorts_3_11_8_en,
    output[1:0] io_VwirePorts_3_11_8_out,
    input [1:0] io_VwirePorts_3_11_7_in,
    input  io_VwirePorts_3_11_7_en,
    output[1:0] io_VwirePorts_3_11_7_out,
    input [1:0] io_VwirePorts_3_11_6_in,
    input  io_VwirePorts_3_11_6_en,
    output[1:0] io_VwirePorts_3_11_6_out,
    input [1:0] io_VwirePorts_3_11_5_in,
    input  io_VwirePorts_3_11_5_en,
    output[1:0] io_VwirePorts_3_11_5_out,
    input [1:0] io_VwirePorts_3_11_4_in,
    input  io_VwirePorts_3_11_4_en,
    output[1:0] io_VwirePorts_3_11_4_out,
    input [1:0] io_VwirePorts_3_11_3_in,
    input  io_VwirePorts_3_11_3_en,
    output[1:0] io_VwirePorts_3_11_3_out,
    input [1:0] io_VwirePorts_3_11_2_in,
    input  io_VwirePorts_3_11_2_en,
    output[1:0] io_VwirePorts_3_11_2_out,
    input [1:0] io_VwirePorts_3_11_1_in,
    input  io_VwirePorts_3_11_1_en,
    output[1:0] io_VwirePorts_3_11_1_out,
    input [1:0] io_VwirePorts_3_11_0_in,
    input  io_VwirePorts_3_11_0_en,
    output[1:0] io_VwirePorts_3_11_0_out,
    input [1:0] io_VwirePorts_3_10_15_in,
    input  io_VwirePorts_3_10_15_en,
    output[1:0] io_VwirePorts_3_10_15_out,
    input [1:0] io_VwirePorts_3_10_14_in,
    input  io_VwirePorts_3_10_14_en,
    output[1:0] io_VwirePorts_3_10_14_out,
    input [1:0] io_VwirePorts_3_10_13_in,
    input  io_VwirePorts_3_10_13_en,
    output[1:0] io_VwirePorts_3_10_13_out,
    input [1:0] io_VwirePorts_3_10_12_in,
    input  io_VwirePorts_3_10_12_en,
    output[1:0] io_VwirePorts_3_10_12_out,
    input [1:0] io_VwirePorts_3_10_11_in,
    input  io_VwirePorts_3_10_11_en,
    output[1:0] io_VwirePorts_3_10_11_out,
    input [1:0] io_VwirePorts_3_10_10_in,
    input  io_VwirePorts_3_10_10_en,
    output[1:0] io_VwirePorts_3_10_10_out,
    input [1:0] io_VwirePorts_3_10_9_in,
    input  io_VwirePorts_3_10_9_en,
    output[1:0] io_VwirePorts_3_10_9_out,
    input [1:0] io_VwirePorts_3_10_8_in,
    input  io_VwirePorts_3_10_8_en,
    output[1:0] io_VwirePorts_3_10_8_out,
    input [1:0] io_VwirePorts_3_10_7_in,
    input  io_VwirePorts_3_10_7_en,
    output[1:0] io_VwirePorts_3_10_7_out,
    input [1:0] io_VwirePorts_3_10_6_in,
    input  io_VwirePorts_3_10_6_en,
    output[1:0] io_VwirePorts_3_10_6_out,
    input [1:0] io_VwirePorts_3_10_5_in,
    input  io_VwirePorts_3_10_5_en,
    output[1:0] io_VwirePorts_3_10_5_out,
    input [1:0] io_VwirePorts_3_10_4_in,
    input  io_VwirePorts_3_10_4_en,
    output[1:0] io_VwirePorts_3_10_4_out,
    input [1:0] io_VwirePorts_3_10_3_in,
    input  io_VwirePorts_3_10_3_en,
    output[1:0] io_VwirePorts_3_10_3_out,
    input [1:0] io_VwirePorts_3_10_2_in,
    input  io_VwirePorts_3_10_2_en,
    output[1:0] io_VwirePorts_3_10_2_out,
    input [1:0] io_VwirePorts_3_10_1_in,
    input  io_VwirePorts_3_10_1_en,
    output[1:0] io_VwirePorts_3_10_1_out,
    input [1:0] io_VwirePorts_3_10_0_in,
    input  io_VwirePorts_3_10_0_en,
    output[1:0] io_VwirePorts_3_10_0_out,
    input [1:0] io_VwirePorts_3_9_15_in,
    input  io_VwirePorts_3_9_15_en,
    output[1:0] io_VwirePorts_3_9_15_out,
    input [1:0] io_VwirePorts_3_9_14_in,
    input  io_VwirePorts_3_9_14_en,
    output[1:0] io_VwirePorts_3_9_14_out,
    input [1:0] io_VwirePorts_3_9_13_in,
    input  io_VwirePorts_3_9_13_en,
    output[1:0] io_VwirePorts_3_9_13_out,
    input [1:0] io_VwirePorts_3_9_12_in,
    input  io_VwirePorts_3_9_12_en,
    output[1:0] io_VwirePorts_3_9_12_out,
    input [1:0] io_VwirePorts_3_9_11_in,
    input  io_VwirePorts_3_9_11_en,
    output[1:0] io_VwirePorts_3_9_11_out,
    input [1:0] io_VwirePorts_3_9_10_in,
    input  io_VwirePorts_3_9_10_en,
    output[1:0] io_VwirePorts_3_9_10_out,
    input [1:0] io_VwirePorts_3_9_9_in,
    input  io_VwirePorts_3_9_9_en,
    output[1:0] io_VwirePorts_3_9_9_out,
    input [1:0] io_VwirePorts_3_9_8_in,
    input  io_VwirePorts_3_9_8_en,
    output[1:0] io_VwirePorts_3_9_8_out,
    input [1:0] io_VwirePorts_3_9_7_in,
    input  io_VwirePorts_3_9_7_en,
    output[1:0] io_VwirePorts_3_9_7_out,
    input [1:0] io_VwirePorts_3_9_6_in,
    input  io_VwirePorts_3_9_6_en,
    output[1:0] io_VwirePorts_3_9_6_out,
    input [1:0] io_VwirePorts_3_9_5_in,
    input  io_VwirePorts_3_9_5_en,
    output[1:0] io_VwirePorts_3_9_5_out,
    input [1:0] io_VwirePorts_3_9_4_in,
    input  io_VwirePorts_3_9_4_en,
    output[1:0] io_VwirePorts_3_9_4_out,
    input [1:0] io_VwirePorts_3_9_3_in,
    input  io_VwirePorts_3_9_3_en,
    output[1:0] io_VwirePorts_3_9_3_out,
    input [1:0] io_VwirePorts_3_9_2_in,
    input  io_VwirePorts_3_9_2_en,
    output[1:0] io_VwirePorts_3_9_2_out,
    input [1:0] io_VwirePorts_3_9_1_in,
    input  io_VwirePorts_3_9_1_en,
    output[1:0] io_VwirePorts_3_9_1_out,
    input [1:0] io_VwirePorts_3_9_0_in,
    input  io_VwirePorts_3_9_0_en,
    output[1:0] io_VwirePorts_3_9_0_out,
    input [1:0] io_VwirePorts_3_8_15_in,
    input  io_VwirePorts_3_8_15_en,
    output[1:0] io_VwirePorts_3_8_15_out,
    input [1:0] io_VwirePorts_3_8_14_in,
    input  io_VwirePorts_3_8_14_en,
    output[1:0] io_VwirePorts_3_8_14_out,
    input [1:0] io_VwirePorts_3_8_13_in,
    input  io_VwirePorts_3_8_13_en,
    output[1:0] io_VwirePorts_3_8_13_out,
    input [1:0] io_VwirePorts_3_8_12_in,
    input  io_VwirePorts_3_8_12_en,
    output[1:0] io_VwirePorts_3_8_12_out,
    input [1:0] io_VwirePorts_3_8_11_in,
    input  io_VwirePorts_3_8_11_en,
    output[1:0] io_VwirePorts_3_8_11_out,
    input [1:0] io_VwirePorts_3_8_10_in,
    input  io_VwirePorts_3_8_10_en,
    output[1:0] io_VwirePorts_3_8_10_out,
    input [1:0] io_VwirePorts_3_8_9_in,
    input  io_VwirePorts_3_8_9_en,
    output[1:0] io_VwirePorts_3_8_9_out,
    input [1:0] io_VwirePorts_3_8_8_in,
    input  io_VwirePorts_3_8_8_en,
    output[1:0] io_VwirePorts_3_8_8_out,
    input [1:0] io_VwirePorts_3_8_7_in,
    input  io_VwirePorts_3_8_7_en,
    output[1:0] io_VwirePorts_3_8_7_out,
    input [1:0] io_VwirePorts_3_8_6_in,
    input  io_VwirePorts_3_8_6_en,
    output[1:0] io_VwirePorts_3_8_6_out,
    input [1:0] io_VwirePorts_3_8_5_in,
    input  io_VwirePorts_3_8_5_en,
    output[1:0] io_VwirePorts_3_8_5_out,
    input [1:0] io_VwirePorts_3_8_4_in,
    input  io_VwirePorts_3_8_4_en,
    output[1:0] io_VwirePorts_3_8_4_out,
    input [1:0] io_VwirePorts_3_8_3_in,
    input  io_VwirePorts_3_8_3_en,
    output[1:0] io_VwirePorts_3_8_3_out,
    input [1:0] io_VwirePorts_3_8_2_in,
    input  io_VwirePorts_3_8_2_en,
    output[1:0] io_VwirePorts_3_8_2_out,
    input [1:0] io_VwirePorts_3_8_1_in,
    input  io_VwirePorts_3_8_1_en,
    output[1:0] io_VwirePorts_3_8_1_out,
    input [1:0] io_VwirePorts_3_8_0_in,
    input  io_VwirePorts_3_8_0_en,
    output[1:0] io_VwirePorts_3_8_0_out,
    input [1:0] io_VwirePorts_3_7_15_in,
    input  io_VwirePorts_3_7_15_en,
    output[1:0] io_VwirePorts_3_7_15_out,
    input [1:0] io_VwirePorts_3_7_14_in,
    input  io_VwirePorts_3_7_14_en,
    output[1:0] io_VwirePorts_3_7_14_out,
    input [1:0] io_VwirePorts_3_7_13_in,
    input  io_VwirePorts_3_7_13_en,
    output[1:0] io_VwirePorts_3_7_13_out,
    input [1:0] io_VwirePorts_3_7_12_in,
    input  io_VwirePorts_3_7_12_en,
    output[1:0] io_VwirePorts_3_7_12_out,
    input [1:0] io_VwirePorts_3_7_11_in,
    input  io_VwirePorts_3_7_11_en,
    output[1:0] io_VwirePorts_3_7_11_out,
    input [1:0] io_VwirePorts_3_7_10_in,
    input  io_VwirePorts_3_7_10_en,
    output[1:0] io_VwirePorts_3_7_10_out,
    input [1:0] io_VwirePorts_3_7_9_in,
    input  io_VwirePorts_3_7_9_en,
    output[1:0] io_VwirePorts_3_7_9_out,
    input [1:0] io_VwirePorts_3_7_8_in,
    input  io_VwirePorts_3_7_8_en,
    output[1:0] io_VwirePorts_3_7_8_out,
    input [1:0] io_VwirePorts_3_7_7_in,
    input  io_VwirePorts_3_7_7_en,
    output[1:0] io_VwirePorts_3_7_7_out,
    input [1:0] io_VwirePorts_3_7_6_in,
    input  io_VwirePorts_3_7_6_en,
    output[1:0] io_VwirePorts_3_7_6_out,
    input [1:0] io_VwirePorts_3_7_5_in,
    input  io_VwirePorts_3_7_5_en,
    output[1:0] io_VwirePorts_3_7_5_out,
    input [1:0] io_VwirePorts_3_7_4_in,
    input  io_VwirePorts_3_7_4_en,
    output[1:0] io_VwirePorts_3_7_4_out,
    input [1:0] io_VwirePorts_3_7_3_in,
    input  io_VwirePorts_3_7_3_en,
    output[1:0] io_VwirePorts_3_7_3_out,
    input [1:0] io_VwirePorts_3_7_2_in,
    input  io_VwirePorts_3_7_2_en,
    output[1:0] io_VwirePorts_3_7_2_out,
    input [1:0] io_VwirePorts_3_7_1_in,
    input  io_VwirePorts_3_7_1_en,
    output[1:0] io_VwirePorts_3_7_1_out,
    input [1:0] io_VwirePorts_3_7_0_in,
    input  io_VwirePorts_3_7_0_en,
    output[1:0] io_VwirePorts_3_7_0_out,
    input [1:0] io_VwirePorts_3_6_15_in,
    input  io_VwirePorts_3_6_15_en,
    output[1:0] io_VwirePorts_3_6_15_out,
    input [1:0] io_VwirePorts_3_6_14_in,
    input  io_VwirePorts_3_6_14_en,
    output[1:0] io_VwirePorts_3_6_14_out,
    input [1:0] io_VwirePorts_3_6_13_in,
    input  io_VwirePorts_3_6_13_en,
    output[1:0] io_VwirePorts_3_6_13_out,
    input [1:0] io_VwirePorts_3_6_12_in,
    input  io_VwirePorts_3_6_12_en,
    output[1:0] io_VwirePorts_3_6_12_out,
    input [1:0] io_VwirePorts_3_6_11_in,
    input  io_VwirePorts_3_6_11_en,
    output[1:0] io_VwirePorts_3_6_11_out,
    input [1:0] io_VwirePorts_3_6_10_in,
    input  io_VwirePorts_3_6_10_en,
    output[1:0] io_VwirePorts_3_6_10_out,
    input [1:0] io_VwirePorts_3_6_9_in,
    input  io_VwirePorts_3_6_9_en,
    output[1:0] io_VwirePorts_3_6_9_out,
    input [1:0] io_VwirePorts_3_6_8_in,
    input  io_VwirePorts_3_6_8_en,
    output[1:0] io_VwirePorts_3_6_8_out,
    input [1:0] io_VwirePorts_3_6_7_in,
    input  io_VwirePorts_3_6_7_en,
    output[1:0] io_VwirePorts_3_6_7_out,
    input [1:0] io_VwirePorts_3_6_6_in,
    input  io_VwirePorts_3_6_6_en,
    output[1:0] io_VwirePorts_3_6_6_out,
    input [1:0] io_VwirePorts_3_6_5_in,
    input  io_VwirePorts_3_6_5_en,
    output[1:0] io_VwirePorts_3_6_5_out,
    input [1:0] io_VwirePorts_3_6_4_in,
    input  io_VwirePorts_3_6_4_en,
    output[1:0] io_VwirePorts_3_6_4_out,
    input [1:0] io_VwirePorts_3_6_3_in,
    input  io_VwirePorts_3_6_3_en,
    output[1:0] io_VwirePorts_3_6_3_out,
    input [1:0] io_VwirePorts_3_6_2_in,
    input  io_VwirePorts_3_6_2_en,
    output[1:0] io_VwirePorts_3_6_2_out,
    input [1:0] io_VwirePorts_3_6_1_in,
    input  io_VwirePorts_3_6_1_en,
    output[1:0] io_VwirePorts_3_6_1_out,
    input [1:0] io_VwirePorts_3_6_0_in,
    input  io_VwirePorts_3_6_0_en,
    output[1:0] io_VwirePorts_3_6_0_out,
    input [1:0] io_VwirePorts_3_5_15_in,
    input  io_VwirePorts_3_5_15_en,
    output[1:0] io_VwirePorts_3_5_15_out,
    input [1:0] io_VwirePorts_3_5_14_in,
    input  io_VwirePorts_3_5_14_en,
    output[1:0] io_VwirePorts_3_5_14_out,
    input [1:0] io_VwirePorts_3_5_13_in,
    input  io_VwirePorts_3_5_13_en,
    output[1:0] io_VwirePorts_3_5_13_out,
    input [1:0] io_VwirePorts_3_5_12_in,
    input  io_VwirePorts_3_5_12_en,
    output[1:0] io_VwirePorts_3_5_12_out,
    input [1:0] io_VwirePorts_3_5_11_in,
    input  io_VwirePorts_3_5_11_en,
    output[1:0] io_VwirePorts_3_5_11_out,
    input [1:0] io_VwirePorts_3_5_10_in,
    input  io_VwirePorts_3_5_10_en,
    output[1:0] io_VwirePorts_3_5_10_out,
    input [1:0] io_VwirePorts_3_5_9_in,
    input  io_VwirePorts_3_5_9_en,
    output[1:0] io_VwirePorts_3_5_9_out,
    input [1:0] io_VwirePorts_3_5_8_in,
    input  io_VwirePorts_3_5_8_en,
    output[1:0] io_VwirePorts_3_5_8_out,
    input [1:0] io_VwirePorts_3_5_7_in,
    input  io_VwirePorts_3_5_7_en,
    output[1:0] io_VwirePorts_3_5_7_out,
    input [1:0] io_VwirePorts_3_5_6_in,
    input  io_VwirePorts_3_5_6_en,
    output[1:0] io_VwirePorts_3_5_6_out,
    input [1:0] io_VwirePorts_3_5_5_in,
    input  io_VwirePorts_3_5_5_en,
    output[1:0] io_VwirePorts_3_5_5_out,
    input [1:0] io_VwirePorts_3_5_4_in,
    input  io_VwirePorts_3_5_4_en,
    output[1:0] io_VwirePorts_3_5_4_out,
    input [1:0] io_VwirePorts_3_5_3_in,
    input  io_VwirePorts_3_5_3_en,
    output[1:0] io_VwirePorts_3_5_3_out,
    input [1:0] io_VwirePorts_3_5_2_in,
    input  io_VwirePorts_3_5_2_en,
    output[1:0] io_VwirePorts_3_5_2_out,
    input [1:0] io_VwirePorts_3_5_1_in,
    input  io_VwirePorts_3_5_1_en,
    output[1:0] io_VwirePorts_3_5_1_out,
    input [1:0] io_VwirePorts_3_5_0_in,
    input  io_VwirePorts_3_5_0_en,
    output[1:0] io_VwirePorts_3_5_0_out,
    input [1:0] io_VwirePorts_3_4_15_in,
    input  io_VwirePorts_3_4_15_en,
    output[1:0] io_VwirePorts_3_4_15_out,
    input [1:0] io_VwirePorts_3_4_14_in,
    input  io_VwirePorts_3_4_14_en,
    output[1:0] io_VwirePorts_3_4_14_out,
    input [1:0] io_VwirePorts_3_4_13_in,
    input  io_VwirePorts_3_4_13_en,
    output[1:0] io_VwirePorts_3_4_13_out,
    input [1:0] io_VwirePorts_3_4_12_in,
    input  io_VwirePorts_3_4_12_en,
    output[1:0] io_VwirePorts_3_4_12_out,
    input [1:0] io_VwirePorts_3_4_11_in,
    input  io_VwirePorts_3_4_11_en,
    output[1:0] io_VwirePorts_3_4_11_out,
    input [1:0] io_VwirePorts_3_4_10_in,
    input  io_VwirePorts_3_4_10_en,
    output[1:0] io_VwirePorts_3_4_10_out,
    input [1:0] io_VwirePorts_3_4_9_in,
    input  io_VwirePorts_3_4_9_en,
    output[1:0] io_VwirePorts_3_4_9_out,
    input [1:0] io_VwirePorts_3_4_8_in,
    input  io_VwirePorts_3_4_8_en,
    output[1:0] io_VwirePorts_3_4_8_out,
    input [1:0] io_VwirePorts_3_4_7_in,
    input  io_VwirePorts_3_4_7_en,
    output[1:0] io_VwirePorts_3_4_7_out,
    input [1:0] io_VwirePorts_3_4_6_in,
    input  io_VwirePorts_3_4_6_en,
    output[1:0] io_VwirePorts_3_4_6_out,
    input [1:0] io_VwirePorts_3_4_5_in,
    input  io_VwirePorts_3_4_5_en,
    output[1:0] io_VwirePorts_3_4_5_out,
    input [1:0] io_VwirePorts_3_4_4_in,
    input  io_VwirePorts_3_4_4_en,
    output[1:0] io_VwirePorts_3_4_4_out,
    input [1:0] io_VwirePorts_3_4_3_in,
    input  io_VwirePorts_3_4_3_en,
    output[1:0] io_VwirePorts_3_4_3_out,
    input [1:0] io_VwirePorts_3_4_2_in,
    input  io_VwirePorts_3_4_2_en,
    output[1:0] io_VwirePorts_3_4_2_out,
    input [1:0] io_VwirePorts_3_4_1_in,
    input  io_VwirePorts_3_4_1_en,
    output[1:0] io_VwirePorts_3_4_1_out,
    input [1:0] io_VwirePorts_3_4_0_in,
    input  io_VwirePorts_3_4_0_en,
    output[1:0] io_VwirePorts_3_4_0_out,
    input [1:0] io_VwirePorts_3_3_15_in,
    input  io_VwirePorts_3_3_15_en,
    output[1:0] io_VwirePorts_3_3_15_out,
    input [1:0] io_VwirePorts_3_3_14_in,
    input  io_VwirePorts_3_3_14_en,
    output[1:0] io_VwirePorts_3_3_14_out,
    input [1:0] io_VwirePorts_3_3_13_in,
    input  io_VwirePorts_3_3_13_en,
    output[1:0] io_VwirePorts_3_3_13_out,
    input [1:0] io_VwirePorts_3_3_12_in,
    input  io_VwirePorts_3_3_12_en,
    output[1:0] io_VwirePorts_3_3_12_out,
    input [1:0] io_VwirePorts_3_3_11_in,
    input  io_VwirePorts_3_3_11_en,
    output[1:0] io_VwirePorts_3_3_11_out,
    input [1:0] io_VwirePorts_3_3_10_in,
    input  io_VwirePorts_3_3_10_en,
    output[1:0] io_VwirePorts_3_3_10_out,
    input [1:0] io_VwirePorts_3_3_9_in,
    input  io_VwirePorts_3_3_9_en,
    output[1:0] io_VwirePorts_3_3_9_out,
    input [1:0] io_VwirePorts_3_3_8_in,
    input  io_VwirePorts_3_3_8_en,
    output[1:0] io_VwirePorts_3_3_8_out,
    input [1:0] io_VwirePorts_3_3_7_in,
    input  io_VwirePorts_3_3_7_en,
    output[1:0] io_VwirePorts_3_3_7_out,
    input [1:0] io_VwirePorts_3_3_6_in,
    input  io_VwirePorts_3_3_6_en,
    output[1:0] io_VwirePorts_3_3_6_out,
    input [1:0] io_VwirePorts_3_3_5_in,
    input  io_VwirePorts_3_3_5_en,
    output[1:0] io_VwirePorts_3_3_5_out,
    input [1:0] io_VwirePorts_3_3_4_in,
    input  io_VwirePorts_3_3_4_en,
    output[1:0] io_VwirePorts_3_3_4_out,
    input [1:0] io_VwirePorts_3_3_3_in,
    input  io_VwirePorts_3_3_3_en,
    output[1:0] io_VwirePorts_3_3_3_out,
    input [1:0] io_VwirePorts_3_3_2_in,
    input  io_VwirePorts_3_3_2_en,
    output[1:0] io_VwirePorts_3_3_2_out,
    input [1:0] io_VwirePorts_3_3_1_in,
    input  io_VwirePorts_3_3_1_en,
    output[1:0] io_VwirePorts_3_3_1_out,
    input [1:0] io_VwirePorts_3_3_0_in,
    input  io_VwirePorts_3_3_0_en,
    output[1:0] io_VwirePorts_3_3_0_out,
    input [1:0] io_VwirePorts_3_2_15_in,
    input  io_VwirePorts_3_2_15_en,
    output[1:0] io_VwirePorts_3_2_15_out,
    input [1:0] io_VwirePorts_3_2_14_in,
    input  io_VwirePorts_3_2_14_en,
    output[1:0] io_VwirePorts_3_2_14_out,
    input [1:0] io_VwirePorts_3_2_13_in,
    input  io_VwirePorts_3_2_13_en,
    output[1:0] io_VwirePorts_3_2_13_out,
    input [1:0] io_VwirePorts_3_2_12_in,
    input  io_VwirePorts_3_2_12_en,
    output[1:0] io_VwirePorts_3_2_12_out,
    input [1:0] io_VwirePorts_3_2_11_in,
    input  io_VwirePorts_3_2_11_en,
    output[1:0] io_VwirePorts_3_2_11_out,
    input [1:0] io_VwirePorts_3_2_10_in,
    input  io_VwirePorts_3_2_10_en,
    output[1:0] io_VwirePorts_3_2_10_out,
    input [1:0] io_VwirePorts_3_2_9_in,
    input  io_VwirePorts_3_2_9_en,
    output[1:0] io_VwirePorts_3_2_9_out,
    input [1:0] io_VwirePorts_3_2_8_in,
    input  io_VwirePorts_3_2_8_en,
    output[1:0] io_VwirePorts_3_2_8_out,
    input [1:0] io_VwirePorts_3_2_7_in,
    input  io_VwirePorts_3_2_7_en,
    output[1:0] io_VwirePorts_3_2_7_out,
    input [1:0] io_VwirePorts_3_2_6_in,
    input  io_VwirePorts_3_2_6_en,
    output[1:0] io_VwirePorts_3_2_6_out,
    input [1:0] io_VwirePorts_3_2_5_in,
    input  io_VwirePorts_3_2_5_en,
    output[1:0] io_VwirePorts_3_2_5_out,
    input [1:0] io_VwirePorts_3_2_4_in,
    input  io_VwirePorts_3_2_4_en,
    output[1:0] io_VwirePorts_3_2_4_out,
    input [1:0] io_VwirePorts_3_2_3_in,
    input  io_VwirePorts_3_2_3_en,
    output[1:0] io_VwirePorts_3_2_3_out,
    input [1:0] io_VwirePorts_3_2_2_in,
    input  io_VwirePorts_3_2_2_en,
    output[1:0] io_VwirePorts_3_2_2_out,
    input [1:0] io_VwirePorts_3_2_1_in,
    input  io_VwirePorts_3_2_1_en,
    output[1:0] io_VwirePorts_3_2_1_out,
    input [1:0] io_VwirePorts_3_2_0_in,
    input  io_VwirePorts_3_2_0_en,
    output[1:0] io_VwirePorts_3_2_0_out,
    input [1:0] io_VwirePorts_3_1_15_in,
    input  io_VwirePorts_3_1_15_en,
    output[1:0] io_VwirePorts_3_1_15_out,
    input [1:0] io_VwirePorts_3_1_14_in,
    input  io_VwirePorts_3_1_14_en,
    output[1:0] io_VwirePorts_3_1_14_out,
    input [1:0] io_VwirePorts_3_1_13_in,
    input  io_VwirePorts_3_1_13_en,
    output[1:0] io_VwirePorts_3_1_13_out,
    input [1:0] io_VwirePorts_3_1_12_in,
    input  io_VwirePorts_3_1_12_en,
    output[1:0] io_VwirePorts_3_1_12_out,
    input [1:0] io_VwirePorts_3_1_11_in,
    input  io_VwirePorts_3_1_11_en,
    output[1:0] io_VwirePorts_3_1_11_out,
    input [1:0] io_VwirePorts_3_1_10_in,
    input  io_VwirePorts_3_1_10_en,
    output[1:0] io_VwirePorts_3_1_10_out,
    input [1:0] io_VwirePorts_3_1_9_in,
    input  io_VwirePorts_3_1_9_en,
    output[1:0] io_VwirePorts_3_1_9_out,
    input [1:0] io_VwirePorts_3_1_8_in,
    input  io_VwirePorts_3_1_8_en,
    output[1:0] io_VwirePorts_3_1_8_out,
    input [1:0] io_VwirePorts_3_1_7_in,
    input  io_VwirePorts_3_1_7_en,
    output[1:0] io_VwirePorts_3_1_7_out,
    input [1:0] io_VwirePorts_3_1_6_in,
    input  io_VwirePorts_3_1_6_en,
    output[1:0] io_VwirePorts_3_1_6_out,
    input [1:0] io_VwirePorts_3_1_5_in,
    input  io_VwirePorts_3_1_5_en,
    output[1:0] io_VwirePorts_3_1_5_out,
    input [1:0] io_VwirePorts_3_1_4_in,
    input  io_VwirePorts_3_1_4_en,
    output[1:0] io_VwirePorts_3_1_4_out,
    input [1:0] io_VwirePorts_3_1_3_in,
    input  io_VwirePorts_3_1_3_en,
    output[1:0] io_VwirePorts_3_1_3_out,
    input [1:0] io_VwirePorts_3_1_2_in,
    input  io_VwirePorts_3_1_2_en,
    output[1:0] io_VwirePorts_3_1_2_out,
    input [1:0] io_VwirePorts_3_1_1_in,
    input  io_VwirePorts_3_1_1_en,
    output[1:0] io_VwirePorts_3_1_1_out,
    input [1:0] io_VwirePorts_3_1_0_in,
    input  io_VwirePorts_3_1_0_en,
    output[1:0] io_VwirePorts_3_1_0_out,
    input [1:0] io_VwirePorts_3_0_15_in,
    input  io_VwirePorts_3_0_15_en,
    output[1:0] io_VwirePorts_3_0_15_out,
    input [1:0] io_VwirePorts_3_0_14_in,
    input  io_VwirePorts_3_0_14_en,
    output[1:0] io_VwirePorts_3_0_14_out,
    input [1:0] io_VwirePorts_3_0_13_in,
    input  io_VwirePorts_3_0_13_en,
    output[1:0] io_VwirePorts_3_0_13_out,
    input [1:0] io_VwirePorts_3_0_12_in,
    input  io_VwirePorts_3_0_12_en,
    output[1:0] io_VwirePorts_3_0_12_out,
    input [1:0] io_VwirePorts_3_0_11_in,
    input  io_VwirePorts_3_0_11_en,
    output[1:0] io_VwirePorts_3_0_11_out,
    input [1:0] io_VwirePorts_3_0_10_in,
    input  io_VwirePorts_3_0_10_en,
    output[1:0] io_VwirePorts_3_0_10_out,
    input [1:0] io_VwirePorts_3_0_9_in,
    input  io_VwirePorts_3_0_9_en,
    output[1:0] io_VwirePorts_3_0_9_out,
    input [1:0] io_VwirePorts_3_0_8_in,
    input  io_VwirePorts_3_0_8_en,
    output[1:0] io_VwirePorts_3_0_8_out,
    input [1:0] io_VwirePorts_3_0_7_in,
    input  io_VwirePorts_3_0_7_en,
    output[1:0] io_VwirePorts_3_0_7_out,
    input [1:0] io_VwirePorts_3_0_6_in,
    input  io_VwirePorts_3_0_6_en,
    output[1:0] io_VwirePorts_3_0_6_out,
    input [1:0] io_VwirePorts_3_0_5_in,
    input  io_VwirePorts_3_0_5_en,
    output[1:0] io_VwirePorts_3_0_5_out,
    input [1:0] io_VwirePorts_3_0_4_in,
    input  io_VwirePorts_3_0_4_en,
    output[1:0] io_VwirePorts_3_0_4_out,
    input [1:0] io_VwirePorts_3_0_3_in,
    input  io_VwirePorts_3_0_3_en,
    output[1:0] io_VwirePorts_3_0_3_out,
    input [1:0] io_VwirePorts_3_0_2_in,
    input  io_VwirePorts_3_0_2_en,
    output[1:0] io_VwirePorts_3_0_2_out,
    input [1:0] io_VwirePorts_3_0_1_in,
    input  io_VwirePorts_3_0_1_en,
    output[1:0] io_VwirePorts_3_0_1_out,
    input [1:0] io_VwirePorts_3_0_0_in,
    input  io_VwirePorts_3_0_0_en,
    output[1:0] io_VwirePorts_3_0_0_out,
    input [1:0] io_VwirePorts_2_22_15_in,
    input  io_VwirePorts_2_22_15_en,
    output[1:0] io_VwirePorts_2_22_15_out,
    input [1:0] io_VwirePorts_2_22_14_in,
    input  io_VwirePorts_2_22_14_en,
    output[1:0] io_VwirePorts_2_22_14_out,
    input [1:0] io_VwirePorts_2_22_13_in,
    input  io_VwirePorts_2_22_13_en,
    output[1:0] io_VwirePorts_2_22_13_out,
    input [1:0] io_VwirePorts_2_22_12_in,
    input  io_VwirePorts_2_22_12_en,
    output[1:0] io_VwirePorts_2_22_12_out,
    input [1:0] io_VwirePorts_2_22_11_in,
    input  io_VwirePorts_2_22_11_en,
    output[1:0] io_VwirePorts_2_22_11_out,
    input [1:0] io_VwirePorts_2_22_10_in,
    input  io_VwirePorts_2_22_10_en,
    output[1:0] io_VwirePorts_2_22_10_out,
    input [1:0] io_VwirePorts_2_22_9_in,
    input  io_VwirePorts_2_22_9_en,
    output[1:0] io_VwirePorts_2_22_9_out,
    input [1:0] io_VwirePorts_2_22_8_in,
    input  io_VwirePorts_2_22_8_en,
    output[1:0] io_VwirePorts_2_22_8_out,
    input [1:0] io_VwirePorts_2_22_7_in,
    input  io_VwirePorts_2_22_7_en,
    output[1:0] io_VwirePorts_2_22_7_out,
    input [1:0] io_VwirePorts_2_22_6_in,
    input  io_VwirePorts_2_22_6_en,
    output[1:0] io_VwirePorts_2_22_6_out,
    input [1:0] io_VwirePorts_2_22_5_in,
    input  io_VwirePorts_2_22_5_en,
    output[1:0] io_VwirePorts_2_22_5_out,
    input [1:0] io_VwirePorts_2_22_4_in,
    input  io_VwirePorts_2_22_4_en,
    output[1:0] io_VwirePorts_2_22_4_out,
    input [1:0] io_VwirePorts_2_22_3_in,
    input  io_VwirePorts_2_22_3_en,
    output[1:0] io_VwirePorts_2_22_3_out,
    input [1:0] io_VwirePorts_2_22_2_in,
    input  io_VwirePorts_2_22_2_en,
    output[1:0] io_VwirePorts_2_22_2_out,
    input [1:0] io_VwirePorts_2_22_1_in,
    input  io_VwirePorts_2_22_1_en,
    output[1:0] io_VwirePorts_2_22_1_out,
    input [1:0] io_VwirePorts_2_22_0_in,
    input  io_VwirePorts_2_22_0_en,
    output[1:0] io_VwirePorts_2_22_0_out,
    input [1:0] io_VwirePorts_2_21_15_in,
    input  io_VwirePorts_2_21_15_en,
    output[1:0] io_VwirePorts_2_21_15_out,
    input [1:0] io_VwirePorts_2_21_14_in,
    input  io_VwirePorts_2_21_14_en,
    output[1:0] io_VwirePorts_2_21_14_out,
    input [1:0] io_VwirePorts_2_21_13_in,
    input  io_VwirePorts_2_21_13_en,
    output[1:0] io_VwirePorts_2_21_13_out,
    input [1:0] io_VwirePorts_2_21_12_in,
    input  io_VwirePorts_2_21_12_en,
    output[1:0] io_VwirePorts_2_21_12_out,
    input [1:0] io_VwirePorts_2_21_11_in,
    input  io_VwirePorts_2_21_11_en,
    output[1:0] io_VwirePorts_2_21_11_out,
    input [1:0] io_VwirePorts_2_21_10_in,
    input  io_VwirePorts_2_21_10_en,
    output[1:0] io_VwirePorts_2_21_10_out,
    input [1:0] io_VwirePorts_2_21_9_in,
    input  io_VwirePorts_2_21_9_en,
    output[1:0] io_VwirePorts_2_21_9_out,
    input [1:0] io_VwirePorts_2_21_8_in,
    input  io_VwirePorts_2_21_8_en,
    output[1:0] io_VwirePorts_2_21_8_out,
    input [1:0] io_VwirePorts_2_21_7_in,
    input  io_VwirePorts_2_21_7_en,
    output[1:0] io_VwirePorts_2_21_7_out,
    input [1:0] io_VwirePorts_2_21_6_in,
    input  io_VwirePorts_2_21_6_en,
    output[1:0] io_VwirePorts_2_21_6_out,
    input [1:0] io_VwirePorts_2_21_5_in,
    input  io_VwirePorts_2_21_5_en,
    output[1:0] io_VwirePorts_2_21_5_out,
    input [1:0] io_VwirePorts_2_21_4_in,
    input  io_VwirePorts_2_21_4_en,
    output[1:0] io_VwirePorts_2_21_4_out,
    input [1:0] io_VwirePorts_2_21_3_in,
    input  io_VwirePorts_2_21_3_en,
    output[1:0] io_VwirePorts_2_21_3_out,
    input [1:0] io_VwirePorts_2_21_2_in,
    input  io_VwirePorts_2_21_2_en,
    output[1:0] io_VwirePorts_2_21_2_out,
    input [1:0] io_VwirePorts_2_21_1_in,
    input  io_VwirePorts_2_21_1_en,
    output[1:0] io_VwirePorts_2_21_1_out,
    input [1:0] io_VwirePorts_2_21_0_in,
    input  io_VwirePorts_2_21_0_en,
    output[1:0] io_VwirePorts_2_21_0_out,
    input [1:0] io_VwirePorts_2_20_15_in,
    input  io_VwirePorts_2_20_15_en,
    output[1:0] io_VwirePorts_2_20_15_out,
    input [1:0] io_VwirePorts_2_20_14_in,
    input  io_VwirePorts_2_20_14_en,
    output[1:0] io_VwirePorts_2_20_14_out,
    input [1:0] io_VwirePorts_2_20_13_in,
    input  io_VwirePorts_2_20_13_en,
    output[1:0] io_VwirePorts_2_20_13_out,
    input [1:0] io_VwirePorts_2_20_12_in,
    input  io_VwirePorts_2_20_12_en,
    output[1:0] io_VwirePorts_2_20_12_out,
    input [1:0] io_VwirePorts_2_20_11_in,
    input  io_VwirePorts_2_20_11_en,
    output[1:0] io_VwirePorts_2_20_11_out,
    input [1:0] io_VwirePorts_2_20_10_in,
    input  io_VwirePorts_2_20_10_en,
    output[1:0] io_VwirePorts_2_20_10_out,
    input [1:0] io_VwirePorts_2_20_9_in,
    input  io_VwirePorts_2_20_9_en,
    output[1:0] io_VwirePorts_2_20_9_out,
    input [1:0] io_VwirePorts_2_20_8_in,
    input  io_VwirePorts_2_20_8_en,
    output[1:0] io_VwirePorts_2_20_8_out,
    input [1:0] io_VwirePorts_2_20_7_in,
    input  io_VwirePorts_2_20_7_en,
    output[1:0] io_VwirePorts_2_20_7_out,
    input [1:0] io_VwirePorts_2_20_6_in,
    input  io_VwirePorts_2_20_6_en,
    output[1:0] io_VwirePorts_2_20_6_out,
    input [1:0] io_VwirePorts_2_20_5_in,
    input  io_VwirePorts_2_20_5_en,
    output[1:0] io_VwirePorts_2_20_5_out,
    input [1:0] io_VwirePorts_2_20_4_in,
    input  io_VwirePorts_2_20_4_en,
    output[1:0] io_VwirePorts_2_20_4_out,
    input [1:0] io_VwirePorts_2_20_3_in,
    input  io_VwirePorts_2_20_3_en,
    output[1:0] io_VwirePorts_2_20_3_out,
    input [1:0] io_VwirePorts_2_20_2_in,
    input  io_VwirePorts_2_20_2_en,
    output[1:0] io_VwirePorts_2_20_2_out,
    input [1:0] io_VwirePorts_2_20_1_in,
    input  io_VwirePorts_2_20_1_en,
    output[1:0] io_VwirePorts_2_20_1_out,
    input [1:0] io_VwirePorts_2_20_0_in,
    input  io_VwirePorts_2_20_0_en,
    output[1:0] io_VwirePorts_2_20_0_out,
    input [1:0] io_VwirePorts_2_19_15_in,
    input  io_VwirePorts_2_19_15_en,
    output[1:0] io_VwirePorts_2_19_15_out,
    input [1:0] io_VwirePorts_2_19_14_in,
    input  io_VwirePorts_2_19_14_en,
    output[1:0] io_VwirePorts_2_19_14_out,
    input [1:0] io_VwirePorts_2_19_13_in,
    input  io_VwirePorts_2_19_13_en,
    output[1:0] io_VwirePorts_2_19_13_out,
    input [1:0] io_VwirePorts_2_19_12_in,
    input  io_VwirePorts_2_19_12_en,
    output[1:0] io_VwirePorts_2_19_12_out,
    input [1:0] io_VwirePorts_2_19_11_in,
    input  io_VwirePorts_2_19_11_en,
    output[1:0] io_VwirePorts_2_19_11_out,
    input [1:0] io_VwirePorts_2_19_10_in,
    input  io_VwirePorts_2_19_10_en,
    output[1:0] io_VwirePorts_2_19_10_out,
    input [1:0] io_VwirePorts_2_19_9_in,
    input  io_VwirePorts_2_19_9_en,
    output[1:0] io_VwirePorts_2_19_9_out,
    input [1:0] io_VwirePorts_2_19_8_in,
    input  io_VwirePorts_2_19_8_en,
    output[1:0] io_VwirePorts_2_19_8_out,
    input [1:0] io_VwirePorts_2_19_7_in,
    input  io_VwirePorts_2_19_7_en,
    output[1:0] io_VwirePorts_2_19_7_out,
    input [1:0] io_VwirePorts_2_19_6_in,
    input  io_VwirePorts_2_19_6_en,
    output[1:0] io_VwirePorts_2_19_6_out,
    input [1:0] io_VwirePorts_2_19_5_in,
    input  io_VwirePorts_2_19_5_en,
    output[1:0] io_VwirePorts_2_19_5_out,
    input [1:0] io_VwirePorts_2_19_4_in,
    input  io_VwirePorts_2_19_4_en,
    output[1:0] io_VwirePorts_2_19_4_out,
    input [1:0] io_VwirePorts_2_19_3_in,
    input  io_VwirePorts_2_19_3_en,
    output[1:0] io_VwirePorts_2_19_3_out,
    input [1:0] io_VwirePorts_2_19_2_in,
    input  io_VwirePorts_2_19_2_en,
    output[1:0] io_VwirePorts_2_19_2_out,
    input [1:0] io_VwirePorts_2_19_1_in,
    input  io_VwirePorts_2_19_1_en,
    output[1:0] io_VwirePorts_2_19_1_out,
    input [1:0] io_VwirePorts_2_19_0_in,
    input  io_VwirePorts_2_19_0_en,
    output[1:0] io_VwirePorts_2_19_0_out,
    input [1:0] io_VwirePorts_2_18_15_in,
    input  io_VwirePorts_2_18_15_en,
    output[1:0] io_VwirePorts_2_18_15_out,
    input [1:0] io_VwirePorts_2_18_14_in,
    input  io_VwirePorts_2_18_14_en,
    output[1:0] io_VwirePorts_2_18_14_out,
    input [1:0] io_VwirePorts_2_18_13_in,
    input  io_VwirePorts_2_18_13_en,
    output[1:0] io_VwirePorts_2_18_13_out,
    input [1:0] io_VwirePorts_2_18_12_in,
    input  io_VwirePorts_2_18_12_en,
    output[1:0] io_VwirePorts_2_18_12_out,
    input [1:0] io_VwirePorts_2_18_11_in,
    input  io_VwirePorts_2_18_11_en,
    output[1:0] io_VwirePorts_2_18_11_out,
    input [1:0] io_VwirePorts_2_18_10_in,
    input  io_VwirePorts_2_18_10_en,
    output[1:0] io_VwirePorts_2_18_10_out,
    input [1:0] io_VwirePorts_2_18_9_in,
    input  io_VwirePorts_2_18_9_en,
    output[1:0] io_VwirePorts_2_18_9_out,
    input [1:0] io_VwirePorts_2_18_8_in,
    input  io_VwirePorts_2_18_8_en,
    output[1:0] io_VwirePorts_2_18_8_out,
    input [1:0] io_VwirePorts_2_18_7_in,
    input  io_VwirePorts_2_18_7_en,
    output[1:0] io_VwirePorts_2_18_7_out,
    input [1:0] io_VwirePorts_2_18_6_in,
    input  io_VwirePorts_2_18_6_en,
    output[1:0] io_VwirePorts_2_18_6_out,
    input [1:0] io_VwirePorts_2_18_5_in,
    input  io_VwirePorts_2_18_5_en,
    output[1:0] io_VwirePorts_2_18_5_out,
    input [1:0] io_VwirePorts_2_18_4_in,
    input  io_VwirePorts_2_18_4_en,
    output[1:0] io_VwirePorts_2_18_4_out,
    input [1:0] io_VwirePorts_2_18_3_in,
    input  io_VwirePorts_2_18_3_en,
    output[1:0] io_VwirePorts_2_18_3_out,
    input [1:0] io_VwirePorts_2_18_2_in,
    input  io_VwirePorts_2_18_2_en,
    output[1:0] io_VwirePorts_2_18_2_out,
    input [1:0] io_VwirePorts_2_18_1_in,
    input  io_VwirePorts_2_18_1_en,
    output[1:0] io_VwirePorts_2_18_1_out,
    input [1:0] io_VwirePorts_2_18_0_in,
    input  io_VwirePorts_2_18_0_en,
    output[1:0] io_VwirePorts_2_18_0_out,
    input [1:0] io_VwirePorts_2_17_15_in,
    input  io_VwirePorts_2_17_15_en,
    output[1:0] io_VwirePorts_2_17_15_out,
    input [1:0] io_VwirePorts_2_17_14_in,
    input  io_VwirePorts_2_17_14_en,
    output[1:0] io_VwirePorts_2_17_14_out,
    input [1:0] io_VwirePorts_2_17_13_in,
    input  io_VwirePorts_2_17_13_en,
    output[1:0] io_VwirePorts_2_17_13_out,
    input [1:0] io_VwirePorts_2_17_12_in,
    input  io_VwirePorts_2_17_12_en,
    output[1:0] io_VwirePorts_2_17_12_out,
    input [1:0] io_VwirePorts_2_17_11_in,
    input  io_VwirePorts_2_17_11_en,
    output[1:0] io_VwirePorts_2_17_11_out,
    input [1:0] io_VwirePorts_2_17_10_in,
    input  io_VwirePorts_2_17_10_en,
    output[1:0] io_VwirePorts_2_17_10_out,
    input [1:0] io_VwirePorts_2_17_9_in,
    input  io_VwirePorts_2_17_9_en,
    output[1:0] io_VwirePorts_2_17_9_out,
    input [1:0] io_VwirePorts_2_17_8_in,
    input  io_VwirePorts_2_17_8_en,
    output[1:0] io_VwirePorts_2_17_8_out,
    input [1:0] io_VwirePorts_2_17_7_in,
    input  io_VwirePorts_2_17_7_en,
    output[1:0] io_VwirePorts_2_17_7_out,
    input [1:0] io_VwirePorts_2_17_6_in,
    input  io_VwirePorts_2_17_6_en,
    output[1:0] io_VwirePorts_2_17_6_out,
    input [1:0] io_VwirePorts_2_17_5_in,
    input  io_VwirePorts_2_17_5_en,
    output[1:0] io_VwirePorts_2_17_5_out,
    input [1:0] io_VwirePorts_2_17_4_in,
    input  io_VwirePorts_2_17_4_en,
    output[1:0] io_VwirePorts_2_17_4_out,
    input [1:0] io_VwirePorts_2_17_3_in,
    input  io_VwirePorts_2_17_3_en,
    output[1:0] io_VwirePorts_2_17_3_out,
    input [1:0] io_VwirePorts_2_17_2_in,
    input  io_VwirePorts_2_17_2_en,
    output[1:0] io_VwirePorts_2_17_2_out,
    input [1:0] io_VwirePorts_2_17_1_in,
    input  io_VwirePorts_2_17_1_en,
    output[1:0] io_VwirePorts_2_17_1_out,
    input [1:0] io_VwirePorts_2_17_0_in,
    input  io_VwirePorts_2_17_0_en,
    output[1:0] io_VwirePorts_2_17_0_out,
    input [1:0] io_VwirePorts_2_16_15_in,
    input  io_VwirePorts_2_16_15_en,
    output[1:0] io_VwirePorts_2_16_15_out,
    input [1:0] io_VwirePorts_2_16_14_in,
    input  io_VwirePorts_2_16_14_en,
    output[1:0] io_VwirePorts_2_16_14_out,
    input [1:0] io_VwirePorts_2_16_13_in,
    input  io_VwirePorts_2_16_13_en,
    output[1:0] io_VwirePorts_2_16_13_out,
    input [1:0] io_VwirePorts_2_16_12_in,
    input  io_VwirePorts_2_16_12_en,
    output[1:0] io_VwirePorts_2_16_12_out,
    input [1:0] io_VwirePorts_2_16_11_in,
    input  io_VwirePorts_2_16_11_en,
    output[1:0] io_VwirePorts_2_16_11_out,
    input [1:0] io_VwirePorts_2_16_10_in,
    input  io_VwirePorts_2_16_10_en,
    output[1:0] io_VwirePorts_2_16_10_out,
    input [1:0] io_VwirePorts_2_16_9_in,
    input  io_VwirePorts_2_16_9_en,
    output[1:0] io_VwirePorts_2_16_9_out,
    input [1:0] io_VwirePorts_2_16_8_in,
    input  io_VwirePorts_2_16_8_en,
    output[1:0] io_VwirePorts_2_16_8_out,
    input [1:0] io_VwirePorts_2_16_7_in,
    input  io_VwirePorts_2_16_7_en,
    output[1:0] io_VwirePorts_2_16_7_out,
    input [1:0] io_VwirePorts_2_16_6_in,
    input  io_VwirePorts_2_16_6_en,
    output[1:0] io_VwirePorts_2_16_6_out,
    input [1:0] io_VwirePorts_2_16_5_in,
    input  io_VwirePorts_2_16_5_en,
    output[1:0] io_VwirePorts_2_16_5_out,
    input [1:0] io_VwirePorts_2_16_4_in,
    input  io_VwirePorts_2_16_4_en,
    output[1:0] io_VwirePorts_2_16_4_out,
    input [1:0] io_VwirePorts_2_16_3_in,
    input  io_VwirePorts_2_16_3_en,
    output[1:0] io_VwirePorts_2_16_3_out,
    input [1:0] io_VwirePorts_2_16_2_in,
    input  io_VwirePorts_2_16_2_en,
    output[1:0] io_VwirePorts_2_16_2_out,
    input [1:0] io_VwirePorts_2_16_1_in,
    input  io_VwirePorts_2_16_1_en,
    output[1:0] io_VwirePorts_2_16_1_out,
    input [1:0] io_VwirePorts_2_16_0_in,
    input  io_VwirePorts_2_16_0_en,
    output[1:0] io_VwirePorts_2_16_0_out,
    input [1:0] io_VwirePorts_2_15_15_in,
    input  io_VwirePorts_2_15_15_en,
    output[1:0] io_VwirePorts_2_15_15_out,
    input [1:0] io_VwirePorts_2_15_14_in,
    input  io_VwirePorts_2_15_14_en,
    output[1:0] io_VwirePorts_2_15_14_out,
    input [1:0] io_VwirePorts_2_15_13_in,
    input  io_VwirePorts_2_15_13_en,
    output[1:0] io_VwirePorts_2_15_13_out,
    input [1:0] io_VwirePorts_2_15_12_in,
    input  io_VwirePorts_2_15_12_en,
    output[1:0] io_VwirePorts_2_15_12_out,
    input [1:0] io_VwirePorts_2_15_11_in,
    input  io_VwirePorts_2_15_11_en,
    output[1:0] io_VwirePorts_2_15_11_out,
    input [1:0] io_VwirePorts_2_15_10_in,
    input  io_VwirePorts_2_15_10_en,
    output[1:0] io_VwirePorts_2_15_10_out,
    input [1:0] io_VwirePorts_2_15_9_in,
    input  io_VwirePorts_2_15_9_en,
    output[1:0] io_VwirePorts_2_15_9_out,
    input [1:0] io_VwirePorts_2_15_8_in,
    input  io_VwirePorts_2_15_8_en,
    output[1:0] io_VwirePorts_2_15_8_out,
    input [1:0] io_VwirePorts_2_15_7_in,
    input  io_VwirePorts_2_15_7_en,
    output[1:0] io_VwirePorts_2_15_7_out,
    input [1:0] io_VwirePorts_2_15_6_in,
    input  io_VwirePorts_2_15_6_en,
    output[1:0] io_VwirePorts_2_15_6_out,
    input [1:0] io_VwirePorts_2_15_5_in,
    input  io_VwirePorts_2_15_5_en,
    output[1:0] io_VwirePorts_2_15_5_out,
    input [1:0] io_VwirePorts_2_15_4_in,
    input  io_VwirePorts_2_15_4_en,
    output[1:0] io_VwirePorts_2_15_4_out,
    input [1:0] io_VwirePorts_2_15_3_in,
    input  io_VwirePorts_2_15_3_en,
    output[1:0] io_VwirePorts_2_15_3_out,
    input [1:0] io_VwirePorts_2_15_2_in,
    input  io_VwirePorts_2_15_2_en,
    output[1:0] io_VwirePorts_2_15_2_out,
    input [1:0] io_VwirePorts_2_15_1_in,
    input  io_VwirePorts_2_15_1_en,
    output[1:0] io_VwirePorts_2_15_1_out,
    input [1:0] io_VwirePorts_2_15_0_in,
    input  io_VwirePorts_2_15_0_en,
    output[1:0] io_VwirePorts_2_15_0_out,
    input [1:0] io_VwirePorts_2_14_15_in,
    input  io_VwirePorts_2_14_15_en,
    output[1:0] io_VwirePorts_2_14_15_out,
    input [1:0] io_VwirePorts_2_14_14_in,
    input  io_VwirePorts_2_14_14_en,
    output[1:0] io_VwirePorts_2_14_14_out,
    input [1:0] io_VwirePorts_2_14_13_in,
    input  io_VwirePorts_2_14_13_en,
    output[1:0] io_VwirePorts_2_14_13_out,
    input [1:0] io_VwirePorts_2_14_12_in,
    input  io_VwirePorts_2_14_12_en,
    output[1:0] io_VwirePorts_2_14_12_out,
    input [1:0] io_VwirePorts_2_14_11_in,
    input  io_VwirePorts_2_14_11_en,
    output[1:0] io_VwirePorts_2_14_11_out,
    input [1:0] io_VwirePorts_2_14_10_in,
    input  io_VwirePorts_2_14_10_en,
    output[1:0] io_VwirePorts_2_14_10_out,
    input [1:0] io_VwirePorts_2_14_9_in,
    input  io_VwirePorts_2_14_9_en,
    output[1:0] io_VwirePorts_2_14_9_out,
    input [1:0] io_VwirePorts_2_14_8_in,
    input  io_VwirePorts_2_14_8_en,
    output[1:0] io_VwirePorts_2_14_8_out,
    input [1:0] io_VwirePorts_2_14_7_in,
    input  io_VwirePorts_2_14_7_en,
    output[1:0] io_VwirePorts_2_14_7_out,
    input [1:0] io_VwirePorts_2_14_6_in,
    input  io_VwirePorts_2_14_6_en,
    output[1:0] io_VwirePorts_2_14_6_out,
    input [1:0] io_VwirePorts_2_14_5_in,
    input  io_VwirePorts_2_14_5_en,
    output[1:0] io_VwirePorts_2_14_5_out,
    input [1:0] io_VwirePorts_2_14_4_in,
    input  io_VwirePorts_2_14_4_en,
    output[1:0] io_VwirePorts_2_14_4_out,
    input [1:0] io_VwirePorts_2_14_3_in,
    input  io_VwirePorts_2_14_3_en,
    output[1:0] io_VwirePorts_2_14_3_out,
    input [1:0] io_VwirePorts_2_14_2_in,
    input  io_VwirePorts_2_14_2_en,
    output[1:0] io_VwirePorts_2_14_2_out,
    input [1:0] io_VwirePorts_2_14_1_in,
    input  io_VwirePorts_2_14_1_en,
    output[1:0] io_VwirePorts_2_14_1_out,
    input [1:0] io_VwirePorts_2_14_0_in,
    input  io_VwirePorts_2_14_0_en,
    output[1:0] io_VwirePorts_2_14_0_out,
    input [1:0] io_VwirePorts_2_13_15_in,
    input  io_VwirePorts_2_13_15_en,
    output[1:0] io_VwirePorts_2_13_15_out,
    input [1:0] io_VwirePorts_2_13_14_in,
    input  io_VwirePorts_2_13_14_en,
    output[1:0] io_VwirePorts_2_13_14_out,
    input [1:0] io_VwirePorts_2_13_13_in,
    input  io_VwirePorts_2_13_13_en,
    output[1:0] io_VwirePorts_2_13_13_out,
    input [1:0] io_VwirePorts_2_13_12_in,
    input  io_VwirePorts_2_13_12_en,
    output[1:0] io_VwirePorts_2_13_12_out,
    input [1:0] io_VwirePorts_2_13_11_in,
    input  io_VwirePorts_2_13_11_en,
    output[1:0] io_VwirePorts_2_13_11_out,
    input [1:0] io_VwirePorts_2_13_10_in,
    input  io_VwirePorts_2_13_10_en,
    output[1:0] io_VwirePorts_2_13_10_out,
    input [1:0] io_VwirePorts_2_13_9_in,
    input  io_VwirePorts_2_13_9_en,
    output[1:0] io_VwirePorts_2_13_9_out,
    input [1:0] io_VwirePorts_2_13_8_in,
    input  io_VwirePorts_2_13_8_en,
    output[1:0] io_VwirePorts_2_13_8_out,
    input [1:0] io_VwirePorts_2_13_7_in,
    input  io_VwirePorts_2_13_7_en,
    output[1:0] io_VwirePorts_2_13_7_out,
    input [1:0] io_VwirePorts_2_13_6_in,
    input  io_VwirePorts_2_13_6_en,
    output[1:0] io_VwirePorts_2_13_6_out,
    input [1:0] io_VwirePorts_2_13_5_in,
    input  io_VwirePorts_2_13_5_en,
    output[1:0] io_VwirePorts_2_13_5_out,
    input [1:0] io_VwirePorts_2_13_4_in,
    input  io_VwirePorts_2_13_4_en,
    output[1:0] io_VwirePorts_2_13_4_out,
    input [1:0] io_VwirePorts_2_13_3_in,
    input  io_VwirePorts_2_13_3_en,
    output[1:0] io_VwirePorts_2_13_3_out,
    input [1:0] io_VwirePorts_2_13_2_in,
    input  io_VwirePorts_2_13_2_en,
    output[1:0] io_VwirePorts_2_13_2_out,
    input [1:0] io_VwirePorts_2_13_1_in,
    input  io_VwirePorts_2_13_1_en,
    output[1:0] io_VwirePorts_2_13_1_out,
    input [1:0] io_VwirePorts_2_13_0_in,
    input  io_VwirePorts_2_13_0_en,
    output[1:0] io_VwirePorts_2_13_0_out,
    input [1:0] io_VwirePorts_2_12_15_in,
    input  io_VwirePorts_2_12_15_en,
    output[1:0] io_VwirePorts_2_12_15_out,
    input [1:0] io_VwirePorts_2_12_14_in,
    input  io_VwirePorts_2_12_14_en,
    output[1:0] io_VwirePorts_2_12_14_out,
    input [1:0] io_VwirePorts_2_12_13_in,
    input  io_VwirePorts_2_12_13_en,
    output[1:0] io_VwirePorts_2_12_13_out,
    input [1:0] io_VwirePorts_2_12_12_in,
    input  io_VwirePorts_2_12_12_en,
    output[1:0] io_VwirePorts_2_12_12_out,
    input [1:0] io_VwirePorts_2_12_11_in,
    input  io_VwirePorts_2_12_11_en,
    output[1:0] io_VwirePorts_2_12_11_out,
    input [1:0] io_VwirePorts_2_12_10_in,
    input  io_VwirePorts_2_12_10_en,
    output[1:0] io_VwirePorts_2_12_10_out,
    input [1:0] io_VwirePorts_2_12_9_in,
    input  io_VwirePorts_2_12_9_en,
    output[1:0] io_VwirePorts_2_12_9_out,
    input [1:0] io_VwirePorts_2_12_8_in,
    input  io_VwirePorts_2_12_8_en,
    output[1:0] io_VwirePorts_2_12_8_out,
    input [1:0] io_VwirePorts_2_12_7_in,
    input  io_VwirePorts_2_12_7_en,
    output[1:0] io_VwirePorts_2_12_7_out,
    input [1:0] io_VwirePorts_2_12_6_in,
    input  io_VwirePorts_2_12_6_en,
    output[1:0] io_VwirePorts_2_12_6_out,
    input [1:0] io_VwirePorts_2_12_5_in,
    input  io_VwirePorts_2_12_5_en,
    output[1:0] io_VwirePorts_2_12_5_out,
    input [1:0] io_VwirePorts_2_12_4_in,
    input  io_VwirePorts_2_12_4_en,
    output[1:0] io_VwirePorts_2_12_4_out,
    input [1:0] io_VwirePorts_2_12_3_in,
    input  io_VwirePorts_2_12_3_en,
    output[1:0] io_VwirePorts_2_12_3_out,
    input [1:0] io_VwirePorts_2_12_2_in,
    input  io_VwirePorts_2_12_2_en,
    output[1:0] io_VwirePorts_2_12_2_out,
    input [1:0] io_VwirePorts_2_12_1_in,
    input  io_VwirePorts_2_12_1_en,
    output[1:0] io_VwirePorts_2_12_1_out,
    input [1:0] io_VwirePorts_2_12_0_in,
    input  io_VwirePorts_2_12_0_en,
    output[1:0] io_VwirePorts_2_12_0_out,
    input [1:0] io_VwirePorts_2_11_15_in,
    input  io_VwirePorts_2_11_15_en,
    output[1:0] io_VwirePorts_2_11_15_out,
    input [1:0] io_VwirePorts_2_11_14_in,
    input  io_VwirePorts_2_11_14_en,
    output[1:0] io_VwirePorts_2_11_14_out,
    input [1:0] io_VwirePorts_2_11_13_in,
    input  io_VwirePorts_2_11_13_en,
    output[1:0] io_VwirePorts_2_11_13_out,
    input [1:0] io_VwirePorts_2_11_12_in,
    input  io_VwirePorts_2_11_12_en,
    output[1:0] io_VwirePorts_2_11_12_out,
    input [1:0] io_VwirePorts_2_11_11_in,
    input  io_VwirePorts_2_11_11_en,
    output[1:0] io_VwirePorts_2_11_11_out,
    input [1:0] io_VwirePorts_2_11_10_in,
    input  io_VwirePorts_2_11_10_en,
    output[1:0] io_VwirePorts_2_11_10_out,
    input [1:0] io_VwirePorts_2_11_9_in,
    input  io_VwirePorts_2_11_9_en,
    output[1:0] io_VwirePorts_2_11_9_out,
    input [1:0] io_VwirePorts_2_11_8_in,
    input  io_VwirePorts_2_11_8_en,
    output[1:0] io_VwirePorts_2_11_8_out,
    input [1:0] io_VwirePorts_2_11_7_in,
    input  io_VwirePorts_2_11_7_en,
    output[1:0] io_VwirePorts_2_11_7_out,
    input [1:0] io_VwirePorts_2_11_6_in,
    input  io_VwirePorts_2_11_6_en,
    output[1:0] io_VwirePorts_2_11_6_out,
    input [1:0] io_VwirePorts_2_11_5_in,
    input  io_VwirePorts_2_11_5_en,
    output[1:0] io_VwirePorts_2_11_5_out,
    input [1:0] io_VwirePorts_2_11_4_in,
    input  io_VwirePorts_2_11_4_en,
    output[1:0] io_VwirePorts_2_11_4_out,
    input [1:0] io_VwirePorts_2_11_3_in,
    input  io_VwirePorts_2_11_3_en,
    output[1:0] io_VwirePorts_2_11_3_out,
    input [1:0] io_VwirePorts_2_11_2_in,
    input  io_VwirePorts_2_11_2_en,
    output[1:0] io_VwirePorts_2_11_2_out,
    input [1:0] io_VwirePorts_2_11_1_in,
    input  io_VwirePorts_2_11_1_en,
    output[1:0] io_VwirePorts_2_11_1_out,
    input [1:0] io_VwirePorts_2_11_0_in,
    input  io_VwirePorts_2_11_0_en,
    output[1:0] io_VwirePorts_2_11_0_out,
    input [1:0] io_VwirePorts_2_10_15_in,
    input  io_VwirePorts_2_10_15_en,
    output[1:0] io_VwirePorts_2_10_15_out,
    input [1:0] io_VwirePorts_2_10_14_in,
    input  io_VwirePorts_2_10_14_en,
    output[1:0] io_VwirePorts_2_10_14_out,
    input [1:0] io_VwirePorts_2_10_13_in,
    input  io_VwirePorts_2_10_13_en,
    output[1:0] io_VwirePorts_2_10_13_out,
    input [1:0] io_VwirePorts_2_10_12_in,
    input  io_VwirePorts_2_10_12_en,
    output[1:0] io_VwirePorts_2_10_12_out,
    input [1:0] io_VwirePorts_2_10_11_in,
    input  io_VwirePorts_2_10_11_en,
    output[1:0] io_VwirePorts_2_10_11_out,
    input [1:0] io_VwirePorts_2_10_10_in,
    input  io_VwirePorts_2_10_10_en,
    output[1:0] io_VwirePorts_2_10_10_out,
    input [1:0] io_VwirePorts_2_10_9_in,
    input  io_VwirePorts_2_10_9_en,
    output[1:0] io_VwirePorts_2_10_9_out,
    input [1:0] io_VwirePorts_2_10_8_in,
    input  io_VwirePorts_2_10_8_en,
    output[1:0] io_VwirePorts_2_10_8_out,
    input [1:0] io_VwirePorts_2_10_7_in,
    input  io_VwirePorts_2_10_7_en,
    output[1:0] io_VwirePorts_2_10_7_out,
    input [1:0] io_VwirePorts_2_10_6_in,
    input  io_VwirePorts_2_10_6_en,
    output[1:0] io_VwirePorts_2_10_6_out,
    input [1:0] io_VwirePorts_2_10_5_in,
    input  io_VwirePorts_2_10_5_en,
    output[1:0] io_VwirePorts_2_10_5_out,
    input [1:0] io_VwirePorts_2_10_4_in,
    input  io_VwirePorts_2_10_4_en,
    output[1:0] io_VwirePorts_2_10_4_out,
    input [1:0] io_VwirePorts_2_10_3_in,
    input  io_VwirePorts_2_10_3_en,
    output[1:0] io_VwirePorts_2_10_3_out,
    input [1:0] io_VwirePorts_2_10_2_in,
    input  io_VwirePorts_2_10_2_en,
    output[1:0] io_VwirePorts_2_10_2_out,
    input [1:0] io_VwirePorts_2_10_1_in,
    input  io_VwirePorts_2_10_1_en,
    output[1:0] io_VwirePorts_2_10_1_out,
    input [1:0] io_VwirePorts_2_10_0_in,
    input  io_VwirePorts_2_10_0_en,
    output[1:0] io_VwirePorts_2_10_0_out,
    input [1:0] io_VwirePorts_2_9_15_in,
    input  io_VwirePorts_2_9_15_en,
    output[1:0] io_VwirePorts_2_9_15_out,
    input [1:0] io_VwirePorts_2_9_14_in,
    input  io_VwirePorts_2_9_14_en,
    output[1:0] io_VwirePorts_2_9_14_out,
    input [1:0] io_VwirePorts_2_9_13_in,
    input  io_VwirePorts_2_9_13_en,
    output[1:0] io_VwirePorts_2_9_13_out,
    input [1:0] io_VwirePorts_2_9_12_in,
    input  io_VwirePorts_2_9_12_en,
    output[1:0] io_VwirePorts_2_9_12_out,
    input [1:0] io_VwirePorts_2_9_11_in,
    input  io_VwirePorts_2_9_11_en,
    output[1:0] io_VwirePorts_2_9_11_out,
    input [1:0] io_VwirePorts_2_9_10_in,
    input  io_VwirePorts_2_9_10_en,
    output[1:0] io_VwirePorts_2_9_10_out,
    input [1:0] io_VwirePorts_2_9_9_in,
    input  io_VwirePorts_2_9_9_en,
    output[1:0] io_VwirePorts_2_9_9_out,
    input [1:0] io_VwirePorts_2_9_8_in,
    input  io_VwirePorts_2_9_8_en,
    output[1:0] io_VwirePorts_2_9_8_out,
    input [1:0] io_VwirePorts_2_9_7_in,
    input  io_VwirePorts_2_9_7_en,
    output[1:0] io_VwirePorts_2_9_7_out,
    input [1:0] io_VwirePorts_2_9_6_in,
    input  io_VwirePorts_2_9_6_en,
    output[1:0] io_VwirePorts_2_9_6_out,
    input [1:0] io_VwirePorts_2_9_5_in,
    input  io_VwirePorts_2_9_5_en,
    output[1:0] io_VwirePorts_2_9_5_out,
    input [1:0] io_VwirePorts_2_9_4_in,
    input  io_VwirePorts_2_9_4_en,
    output[1:0] io_VwirePorts_2_9_4_out,
    input [1:0] io_VwirePorts_2_9_3_in,
    input  io_VwirePorts_2_9_3_en,
    output[1:0] io_VwirePorts_2_9_3_out,
    input [1:0] io_VwirePorts_2_9_2_in,
    input  io_VwirePorts_2_9_2_en,
    output[1:0] io_VwirePorts_2_9_2_out,
    input [1:0] io_VwirePorts_2_9_1_in,
    input  io_VwirePorts_2_9_1_en,
    output[1:0] io_VwirePorts_2_9_1_out,
    input [1:0] io_VwirePorts_2_9_0_in,
    input  io_VwirePorts_2_9_0_en,
    output[1:0] io_VwirePorts_2_9_0_out,
    input [1:0] io_VwirePorts_2_8_15_in,
    input  io_VwirePorts_2_8_15_en,
    output[1:0] io_VwirePorts_2_8_15_out,
    input [1:0] io_VwirePorts_2_8_14_in,
    input  io_VwirePorts_2_8_14_en,
    output[1:0] io_VwirePorts_2_8_14_out,
    input [1:0] io_VwirePorts_2_8_13_in,
    input  io_VwirePorts_2_8_13_en,
    output[1:0] io_VwirePorts_2_8_13_out,
    input [1:0] io_VwirePorts_2_8_12_in,
    input  io_VwirePorts_2_8_12_en,
    output[1:0] io_VwirePorts_2_8_12_out,
    input [1:0] io_VwirePorts_2_8_11_in,
    input  io_VwirePorts_2_8_11_en,
    output[1:0] io_VwirePorts_2_8_11_out,
    input [1:0] io_VwirePorts_2_8_10_in,
    input  io_VwirePorts_2_8_10_en,
    output[1:0] io_VwirePorts_2_8_10_out,
    input [1:0] io_VwirePorts_2_8_9_in,
    input  io_VwirePorts_2_8_9_en,
    output[1:0] io_VwirePorts_2_8_9_out,
    input [1:0] io_VwirePorts_2_8_8_in,
    input  io_VwirePorts_2_8_8_en,
    output[1:0] io_VwirePorts_2_8_8_out,
    input [1:0] io_VwirePorts_2_8_7_in,
    input  io_VwirePorts_2_8_7_en,
    output[1:0] io_VwirePorts_2_8_7_out,
    input [1:0] io_VwirePorts_2_8_6_in,
    input  io_VwirePorts_2_8_6_en,
    output[1:0] io_VwirePorts_2_8_6_out,
    input [1:0] io_VwirePorts_2_8_5_in,
    input  io_VwirePorts_2_8_5_en,
    output[1:0] io_VwirePorts_2_8_5_out,
    input [1:0] io_VwirePorts_2_8_4_in,
    input  io_VwirePorts_2_8_4_en,
    output[1:0] io_VwirePorts_2_8_4_out,
    input [1:0] io_VwirePorts_2_8_3_in,
    input  io_VwirePorts_2_8_3_en,
    output[1:0] io_VwirePorts_2_8_3_out,
    input [1:0] io_VwirePorts_2_8_2_in,
    input  io_VwirePorts_2_8_2_en,
    output[1:0] io_VwirePorts_2_8_2_out,
    input [1:0] io_VwirePorts_2_8_1_in,
    input  io_VwirePorts_2_8_1_en,
    output[1:0] io_VwirePorts_2_8_1_out,
    input [1:0] io_VwirePorts_2_8_0_in,
    input  io_VwirePorts_2_8_0_en,
    output[1:0] io_VwirePorts_2_8_0_out,
    input [1:0] io_VwirePorts_2_7_15_in,
    input  io_VwirePorts_2_7_15_en,
    output[1:0] io_VwirePorts_2_7_15_out,
    input [1:0] io_VwirePorts_2_7_14_in,
    input  io_VwirePorts_2_7_14_en,
    output[1:0] io_VwirePorts_2_7_14_out,
    input [1:0] io_VwirePorts_2_7_13_in,
    input  io_VwirePorts_2_7_13_en,
    output[1:0] io_VwirePorts_2_7_13_out,
    input [1:0] io_VwirePorts_2_7_12_in,
    input  io_VwirePorts_2_7_12_en,
    output[1:0] io_VwirePorts_2_7_12_out,
    input [1:0] io_VwirePorts_2_7_11_in,
    input  io_VwirePorts_2_7_11_en,
    output[1:0] io_VwirePorts_2_7_11_out,
    input [1:0] io_VwirePorts_2_7_10_in,
    input  io_VwirePorts_2_7_10_en,
    output[1:0] io_VwirePorts_2_7_10_out,
    input [1:0] io_VwirePorts_2_7_9_in,
    input  io_VwirePorts_2_7_9_en,
    output[1:0] io_VwirePorts_2_7_9_out,
    input [1:0] io_VwirePorts_2_7_8_in,
    input  io_VwirePorts_2_7_8_en,
    output[1:0] io_VwirePorts_2_7_8_out,
    input [1:0] io_VwirePorts_2_7_7_in,
    input  io_VwirePorts_2_7_7_en,
    output[1:0] io_VwirePorts_2_7_7_out,
    input [1:0] io_VwirePorts_2_7_6_in,
    input  io_VwirePorts_2_7_6_en,
    output[1:0] io_VwirePorts_2_7_6_out,
    input [1:0] io_VwirePorts_2_7_5_in,
    input  io_VwirePorts_2_7_5_en,
    output[1:0] io_VwirePorts_2_7_5_out,
    input [1:0] io_VwirePorts_2_7_4_in,
    input  io_VwirePorts_2_7_4_en,
    output[1:0] io_VwirePorts_2_7_4_out,
    input [1:0] io_VwirePorts_2_7_3_in,
    input  io_VwirePorts_2_7_3_en,
    output[1:0] io_VwirePorts_2_7_3_out,
    input [1:0] io_VwirePorts_2_7_2_in,
    input  io_VwirePorts_2_7_2_en,
    output[1:0] io_VwirePorts_2_7_2_out,
    input [1:0] io_VwirePorts_2_7_1_in,
    input  io_VwirePorts_2_7_1_en,
    output[1:0] io_VwirePorts_2_7_1_out,
    input [1:0] io_VwirePorts_2_7_0_in,
    input  io_VwirePorts_2_7_0_en,
    output[1:0] io_VwirePorts_2_7_0_out,
    input [1:0] io_VwirePorts_2_6_15_in,
    input  io_VwirePorts_2_6_15_en,
    output[1:0] io_VwirePorts_2_6_15_out,
    input [1:0] io_VwirePorts_2_6_14_in,
    input  io_VwirePorts_2_6_14_en,
    output[1:0] io_VwirePorts_2_6_14_out,
    input [1:0] io_VwirePorts_2_6_13_in,
    input  io_VwirePorts_2_6_13_en,
    output[1:0] io_VwirePorts_2_6_13_out,
    input [1:0] io_VwirePorts_2_6_12_in,
    input  io_VwirePorts_2_6_12_en,
    output[1:0] io_VwirePorts_2_6_12_out,
    input [1:0] io_VwirePorts_2_6_11_in,
    input  io_VwirePorts_2_6_11_en,
    output[1:0] io_VwirePorts_2_6_11_out,
    input [1:0] io_VwirePorts_2_6_10_in,
    input  io_VwirePorts_2_6_10_en,
    output[1:0] io_VwirePorts_2_6_10_out,
    input [1:0] io_VwirePorts_2_6_9_in,
    input  io_VwirePorts_2_6_9_en,
    output[1:0] io_VwirePorts_2_6_9_out,
    input [1:0] io_VwirePorts_2_6_8_in,
    input  io_VwirePorts_2_6_8_en,
    output[1:0] io_VwirePorts_2_6_8_out,
    input [1:0] io_VwirePorts_2_6_7_in,
    input  io_VwirePorts_2_6_7_en,
    output[1:0] io_VwirePorts_2_6_7_out,
    input [1:0] io_VwirePorts_2_6_6_in,
    input  io_VwirePorts_2_6_6_en,
    output[1:0] io_VwirePorts_2_6_6_out,
    input [1:0] io_VwirePorts_2_6_5_in,
    input  io_VwirePorts_2_6_5_en,
    output[1:0] io_VwirePorts_2_6_5_out,
    input [1:0] io_VwirePorts_2_6_4_in,
    input  io_VwirePorts_2_6_4_en,
    output[1:0] io_VwirePorts_2_6_4_out,
    input [1:0] io_VwirePorts_2_6_3_in,
    input  io_VwirePorts_2_6_3_en,
    output[1:0] io_VwirePorts_2_6_3_out,
    input [1:0] io_VwirePorts_2_6_2_in,
    input  io_VwirePorts_2_6_2_en,
    output[1:0] io_VwirePorts_2_6_2_out,
    input [1:0] io_VwirePorts_2_6_1_in,
    input  io_VwirePorts_2_6_1_en,
    output[1:0] io_VwirePorts_2_6_1_out,
    input [1:0] io_VwirePorts_2_6_0_in,
    input  io_VwirePorts_2_6_0_en,
    output[1:0] io_VwirePorts_2_6_0_out,
    input [1:0] io_VwirePorts_2_5_15_in,
    input  io_VwirePorts_2_5_15_en,
    output[1:0] io_VwirePorts_2_5_15_out,
    input [1:0] io_VwirePorts_2_5_14_in,
    input  io_VwirePorts_2_5_14_en,
    output[1:0] io_VwirePorts_2_5_14_out,
    input [1:0] io_VwirePorts_2_5_13_in,
    input  io_VwirePorts_2_5_13_en,
    output[1:0] io_VwirePorts_2_5_13_out,
    input [1:0] io_VwirePorts_2_5_12_in,
    input  io_VwirePorts_2_5_12_en,
    output[1:0] io_VwirePorts_2_5_12_out,
    input [1:0] io_VwirePorts_2_5_11_in,
    input  io_VwirePorts_2_5_11_en,
    output[1:0] io_VwirePorts_2_5_11_out,
    input [1:0] io_VwirePorts_2_5_10_in,
    input  io_VwirePorts_2_5_10_en,
    output[1:0] io_VwirePorts_2_5_10_out,
    input [1:0] io_VwirePorts_2_5_9_in,
    input  io_VwirePorts_2_5_9_en,
    output[1:0] io_VwirePorts_2_5_9_out,
    input [1:0] io_VwirePorts_2_5_8_in,
    input  io_VwirePorts_2_5_8_en,
    output[1:0] io_VwirePorts_2_5_8_out,
    input [1:0] io_VwirePorts_2_5_7_in,
    input  io_VwirePorts_2_5_7_en,
    output[1:0] io_VwirePorts_2_5_7_out,
    input [1:0] io_VwirePorts_2_5_6_in,
    input  io_VwirePorts_2_5_6_en,
    output[1:0] io_VwirePorts_2_5_6_out,
    input [1:0] io_VwirePorts_2_5_5_in,
    input  io_VwirePorts_2_5_5_en,
    output[1:0] io_VwirePorts_2_5_5_out,
    input [1:0] io_VwirePorts_2_5_4_in,
    input  io_VwirePorts_2_5_4_en,
    output[1:0] io_VwirePorts_2_5_4_out,
    input [1:0] io_VwirePorts_2_5_3_in,
    input  io_VwirePorts_2_5_3_en,
    output[1:0] io_VwirePorts_2_5_3_out,
    input [1:0] io_VwirePorts_2_5_2_in,
    input  io_VwirePorts_2_5_2_en,
    output[1:0] io_VwirePorts_2_5_2_out,
    input [1:0] io_VwirePorts_2_5_1_in,
    input  io_VwirePorts_2_5_1_en,
    output[1:0] io_VwirePorts_2_5_1_out,
    input [1:0] io_VwirePorts_2_5_0_in,
    input  io_VwirePorts_2_5_0_en,
    output[1:0] io_VwirePorts_2_5_0_out,
    input [1:0] io_VwirePorts_2_4_15_in,
    input  io_VwirePorts_2_4_15_en,
    output[1:0] io_VwirePorts_2_4_15_out,
    input [1:0] io_VwirePorts_2_4_14_in,
    input  io_VwirePorts_2_4_14_en,
    output[1:0] io_VwirePorts_2_4_14_out,
    input [1:0] io_VwirePorts_2_4_13_in,
    input  io_VwirePorts_2_4_13_en,
    output[1:0] io_VwirePorts_2_4_13_out,
    input [1:0] io_VwirePorts_2_4_12_in,
    input  io_VwirePorts_2_4_12_en,
    output[1:0] io_VwirePorts_2_4_12_out,
    input [1:0] io_VwirePorts_2_4_11_in,
    input  io_VwirePorts_2_4_11_en,
    output[1:0] io_VwirePorts_2_4_11_out,
    input [1:0] io_VwirePorts_2_4_10_in,
    input  io_VwirePorts_2_4_10_en,
    output[1:0] io_VwirePorts_2_4_10_out,
    input [1:0] io_VwirePorts_2_4_9_in,
    input  io_VwirePorts_2_4_9_en,
    output[1:0] io_VwirePorts_2_4_9_out,
    input [1:0] io_VwirePorts_2_4_8_in,
    input  io_VwirePorts_2_4_8_en,
    output[1:0] io_VwirePorts_2_4_8_out,
    input [1:0] io_VwirePorts_2_4_7_in,
    input  io_VwirePorts_2_4_7_en,
    output[1:0] io_VwirePorts_2_4_7_out,
    input [1:0] io_VwirePorts_2_4_6_in,
    input  io_VwirePorts_2_4_6_en,
    output[1:0] io_VwirePorts_2_4_6_out,
    input [1:0] io_VwirePorts_2_4_5_in,
    input  io_VwirePorts_2_4_5_en,
    output[1:0] io_VwirePorts_2_4_5_out,
    input [1:0] io_VwirePorts_2_4_4_in,
    input  io_VwirePorts_2_4_4_en,
    output[1:0] io_VwirePorts_2_4_4_out,
    input [1:0] io_VwirePorts_2_4_3_in,
    input  io_VwirePorts_2_4_3_en,
    output[1:0] io_VwirePorts_2_4_3_out,
    input [1:0] io_VwirePorts_2_4_2_in,
    input  io_VwirePorts_2_4_2_en,
    output[1:0] io_VwirePorts_2_4_2_out,
    input [1:0] io_VwirePorts_2_4_1_in,
    input  io_VwirePorts_2_4_1_en,
    output[1:0] io_VwirePorts_2_4_1_out,
    input [1:0] io_VwirePorts_2_4_0_in,
    input  io_VwirePorts_2_4_0_en,
    output[1:0] io_VwirePorts_2_4_0_out,
    input [1:0] io_VwirePorts_2_3_15_in,
    input  io_VwirePorts_2_3_15_en,
    output[1:0] io_VwirePorts_2_3_15_out,
    input [1:0] io_VwirePorts_2_3_14_in,
    input  io_VwirePorts_2_3_14_en,
    output[1:0] io_VwirePorts_2_3_14_out,
    input [1:0] io_VwirePorts_2_3_13_in,
    input  io_VwirePorts_2_3_13_en,
    output[1:0] io_VwirePorts_2_3_13_out,
    input [1:0] io_VwirePorts_2_3_12_in,
    input  io_VwirePorts_2_3_12_en,
    output[1:0] io_VwirePorts_2_3_12_out,
    input [1:0] io_VwirePorts_2_3_11_in,
    input  io_VwirePorts_2_3_11_en,
    output[1:0] io_VwirePorts_2_3_11_out,
    input [1:0] io_VwirePorts_2_3_10_in,
    input  io_VwirePorts_2_3_10_en,
    output[1:0] io_VwirePorts_2_3_10_out,
    input [1:0] io_VwirePorts_2_3_9_in,
    input  io_VwirePorts_2_3_9_en,
    output[1:0] io_VwirePorts_2_3_9_out,
    input [1:0] io_VwirePorts_2_3_8_in,
    input  io_VwirePorts_2_3_8_en,
    output[1:0] io_VwirePorts_2_3_8_out,
    input [1:0] io_VwirePorts_2_3_7_in,
    input  io_VwirePorts_2_3_7_en,
    output[1:0] io_VwirePorts_2_3_7_out,
    input [1:0] io_VwirePorts_2_3_6_in,
    input  io_VwirePorts_2_3_6_en,
    output[1:0] io_VwirePorts_2_3_6_out,
    input [1:0] io_VwirePorts_2_3_5_in,
    input  io_VwirePorts_2_3_5_en,
    output[1:0] io_VwirePorts_2_3_5_out,
    input [1:0] io_VwirePorts_2_3_4_in,
    input  io_VwirePorts_2_3_4_en,
    output[1:0] io_VwirePorts_2_3_4_out,
    input [1:0] io_VwirePorts_2_3_3_in,
    input  io_VwirePorts_2_3_3_en,
    output[1:0] io_VwirePorts_2_3_3_out,
    input [1:0] io_VwirePorts_2_3_2_in,
    input  io_VwirePorts_2_3_2_en,
    output[1:0] io_VwirePorts_2_3_2_out,
    input [1:0] io_VwirePorts_2_3_1_in,
    input  io_VwirePorts_2_3_1_en,
    output[1:0] io_VwirePorts_2_3_1_out,
    input [1:0] io_VwirePorts_2_3_0_in,
    input  io_VwirePorts_2_3_0_en,
    output[1:0] io_VwirePorts_2_3_0_out,
    input [1:0] io_VwirePorts_2_2_15_in,
    input  io_VwirePorts_2_2_15_en,
    output[1:0] io_VwirePorts_2_2_15_out,
    input [1:0] io_VwirePorts_2_2_14_in,
    input  io_VwirePorts_2_2_14_en,
    output[1:0] io_VwirePorts_2_2_14_out,
    input [1:0] io_VwirePorts_2_2_13_in,
    input  io_VwirePorts_2_2_13_en,
    output[1:0] io_VwirePorts_2_2_13_out,
    input [1:0] io_VwirePorts_2_2_12_in,
    input  io_VwirePorts_2_2_12_en,
    output[1:0] io_VwirePorts_2_2_12_out,
    input [1:0] io_VwirePorts_2_2_11_in,
    input  io_VwirePorts_2_2_11_en,
    output[1:0] io_VwirePorts_2_2_11_out,
    input [1:0] io_VwirePorts_2_2_10_in,
    input  io_VwirePorts_2_2_10_en,
    output[1:0] io_VwirePorts_2_2_10_out,
    input [1:0] io_VwirePorts_2_2_9_in,
    input  io_VwirePorts_2_2_9_en,
    output[1:0] io_VwirePorts_2_2_9_out,
    input [1:0] io_VwirePorts_2_2_8_in,
    input  io_VwirePorts_2_2_8_en,
    output[1:0] io_VwirePorts_2_2_8_out,
    input [1:0] io_VwirePorts_2_2_7_in,
    input  io_VwirePorts_2_2_7_en,
    output[1:0] io_VwirePorts_2_2_7_out,
    input [1:0] io_VwirePorts_2_2_6_in,
    input  io_VwirePorts_2_2_6_en,
    output[1:0] io_VwirePorts_2_2_6_out,
    input [1:0] io_VwirePorts_2_2_5_in,
    input  io_VwirePorts_2_2_5_en,
    output[1:0] io_VwirePorts_2_2_5_out,
    input [1:0] io_VwirePorts_2_2_4_in,
    input  io_VwirePorts_2_2_4_en,
    output[1:0] io_VwirePorts_2_2_4_out,
    input [1:0] io_VwirePorts_2_2_3_in,
    input  io_VwirePorts_2_2_3_en,
    output[1:0] io_VwirePorts_2_2_3_out,
    input [1:0] io_VwirePorts_2_2_2_in,
    input  io_VwirePorts_2_2_2_en,
    output[1:0] io_VwirePorts_2_2_2_out,
    input [1:0] io_VwirePorts_2_2_1_in,
    input  io_VwirePorts_2_2_1_en,
    output[1:0] io_VwirePorts_2_2_1_out,
    input [1:0] io_VwirePorts_2_2_0_in,
    input  io_VwirePorts_2_2_0_en,
    output[1:0] io_VwirePorts_2_2_0_out,
    input [1:0] io_VwirePorts_2_1_15_in,
    input  io_VwirePorts_2_1_15_en,
    output[1:0] io_VwirePorts_2_1_15_out,
    input [1:0] io_VwirePorts_2_1_14_in,
    input  io_VwirePorts_2_1_14_en,
    output[1:0] io_VwirePorts_2_1_14_out,
    input [1:0] io_VwirePorts_2_1_13_in,
    input  io_VwirePorts_2_1_13_en,
    output[1:0] io_VwirePorts_2_1_13_out,
    input [1:0] io_VwirePorts_2_1_12_in,
    input  io_VwirePorts_2_1_12_en,
    output[1:0] io_VwirePorts_2_1_12_out,
    input [1:0] io_VwirePorts_2_1_11_in,
    input  io_VwirePorts_2_1_11_en,
    output[1:0] io_VwirePorts_2_1_11_out,
    input [1:0] io_VwirePorts_2_1_10_in,
    input  io_VwirePorts_2_1_10_en,
    output[1:0] io_VwirePorts_2_1_10_out,
    input [1:0] io_VwirePorts_2_1_9_in,
    input  io_VwirePorts_2_1_9_en,
    output[1:0] io_VwirePorts_2_1_9_out,
    input [1:0] io_VwirePorts_2_1_8_in,
    input  io_VwirePorts_2_1_8_en,
    output[1:0] io_VwirePorts_2_1_8_out,
    input [1:0] io_VwirePorts_2_1_7_in,
    input  io_VwirePorts_2_1_7_en,
    output[1:0] io_VwirePorts_2_1_7_out,
    input [1:0] io_VwirePorts_2_1_6_in,
    input  io_VwirePorts_2_1_6_en,
    output[1:0] io_VwirePorts_2_1_6_out,
    input [1:0] io_VwirePorts_2_1_5_in,
    input  io_VwirePorts_2_1_5_en,
    output[1:0] io_VwirePorts_2_1_5_out,
    input [1:0] io_VwirePorts_2_1_4_in,
    input  io_VwirePorts_2_1_4_en,
    output[1:0] io_VwirePorts_2_1_4_out,
    input [1:0] io_VwirePorts_2_1_3_in,
    input  io_VwirePorts_2_1_3_en,
    output[1:0] io_VwirePorts_2_1_3_out,
    input [1:0] io_VwirePorts_2_1_2_in,
    input  io_VwirePorts_2_1_2_en,
    output[1:0] io_VwirePorts_2_1_2_out,
    input [1:0] io_VwirePorts_2_1_1_in,
    input  io_VwirePorts_2_1_1_en,
    output[1:0] io_VwirePorts_2_1_1_out,
    input [1:0] io_VwirePorts_2_1_0_in,
    input  io_VwirePorts_2_1_0_en,
    output[1:0] io_VwirePorts_2_1_0_out,
    input [1:0] io_VwirePorts_2_0_15_in,
    input  io_VwirePorts_2_0_15_en,
    output[1:0] io_VwirePorts_2_0_15_out,
    input [1:0] io_VwirePorts_2_0_14_in,
    input  io_VwirePorts_2_0_14_en,
    output[1:0] io_VwirePorts_2_0_14_out,
    input [1:0] io_VwirePorts_2_0_13_in,
    input  io_VwirePorts_2_0_13_en,
    output[1:0] io_VwirePorts_2_0_13_out,
    input [1:0] io_VwirePorts_2_0_12_in,
    input  io_VwirePorts_2_0_12_en,
    output[1:0] io_VwirePorts_2_0_12_out,
    input [1:0] io_VwirePorts_2_0_11_in,
    input  io_VwirePorts_2_0_11_en,
    output[1:0] io_VwirePorts_2_0_11_out,
    input [1:0] io_VwirePorts_2_0_10_in,
    input  io_VwirePorts_2_0_10_en,
    output[1:0] io_VwirePorts_2_0_10_out,
    input [1:0] io_VwirePorts_2_0_9_in,
    input  io_VwirePorts_2_0_9_en,
    output[1:0] io_VwirePorts_2_0_9_out,
    input [1:0] io_VwirePorts_2_0_8_in,
    input  io_VwirePorts_2_0_8_en,
    output[1:0] io_VwirePorts_2_0_8_out,
    input [1:0] io_VwirePorts_2_0_7_in,
    input  io_VwirePorts_2_0_7_en,
    output[1:0] io_VwirePorts_2_0_7_out,
    input [1:0] io_VwirePorts_2_0_6_in,
    input  io_VwirePorts_2_0_6_en,
    output[1:0] io_VwirePorts_2_0_6_out,
    input [1:0] io_VwirePorts_2_0_5_in,
    input  io_VwirePorts_2_0_5_en,
    output[1:0] io_VwirePorts_2_0_5_out,
    input [1:0] io_VwirePorts_2_0_4_in,
    input  io_VwirePorts_2_0_4_en,
    output[1:0] io_VwirePorts_2_0_4_out,
    input [1:0] io_VwirePorts_2_0_3_in,
    input  io_VwirePorts_2_0_3_en,
    output[1:0] io_VwirePorts_2_0_3_out,
    input [1:0] io_VwirePorts_2_0_2_in,
    input  io_VwirePorts_2_0_2_en,
    output[1:0] io_VwirePorts_2_0_2_out,
    input [1:0] io_VwirePorts_2_0_1_in,
    input  io_VwirePorts_2_0_1_en,
    output[1:0] io_VwirePorts_2_0_1_out,
    input [1:0] io_VwirePorts_2_0_0_in,
    input  io_VwirePorts_2_0_0_en,
    output[1:0] io_VwirePorts_2_0_0_out,
    input [1:0] io_VwirePorts_1_22_15_in,
    input  io_VwirePorts_1_22_15_en,
    output[1:0] io_VwirePorts_1_22_15_out,
    input [1:0] io_VwirePorts_1_22_14_in,
    input  io_VwirePorts_1_22_14_en,
    output[1:0] io_VwirePorts_1_22_14_out,
    input [1:0] io_VwirePorts_1_22_13_in,
    input  io_VwirePorts_1_22_13_en,
    output[1:0] io_VwirePorts_1_22_13_out,
    input [1:0] io_VwirePorts_1_22_12_in,
    input  io_VwirePorts_1_22_12_en,
    output[1:0] io_VwirePorts_1_22_12_out,
    input [1:0] io_VwirePorts_1_22_11_in,
    input  io_VwirePorts_1_22_11_en,
    output[1:0] io_VwirePorts_1_22_11_out,
    input [1:0] io_VwirePorts_1_22_10_in,
    input  io_VwirePorts_1_22_10_en,
    output[1:0] io_VwirePorts_1_22_10_out,
    input [1:0] io_VwirePorts_1_22_9_in,
    input  io_VwirePorts_1_22_9_en,
    output[1:0] io_VwirePorts_1_22_9_out,
    input [1:0] io_VwirePorts_1_22_8_in,
    input  io_VwirePorts_1_22_8_en,
    output[1:0] io_VwirePorts_1_22_8_out,
    input [1:0] io_VwirePorts_1_22_7_in,
    input  io_VwirePorts_1_22_7_en,
    output[1:0] io_VwirePorts_1_22_7_out,
    input [1:0] io_VwirePorts_1_22_6_in,
    input  io_VwirePorts_1_22_6_en,
    output[1:0] io_VwirePorts_1_22_6_out,
    input [1:0] io_VwirePorts_1_22_5_in,
    input  io_VwirePorts_1_22_5_en,
    output[1:0] io_VwirePorts_1_22_5_out,
    input [1:0] io_VwirePorts_1_22_4_in,
    input  io_VwirePorts_1_22_4_en,
    output[1:0] io_VwirePorts_1_22_4_out,
    input [1:0] io_VwirePorts_1_22_3_in,
    input  io_VwirePorts_1_22_3_en,
    output[1:0] io_VwirePorts_1_22_3_out,
    input [1:0] io_VwirePorts_1_22_2_in,
    input  io_VwirePorts_1_22_2_en,
    output[1:0] io_VwirePorts_1_22_2_out,
    input [1:0] io_VwirePorts_1_22_1_in,
    input  io_VwirePorts_1_22_1_en,
    output[1:0] io_VwirePorts_1_22_1_out,
    input [1:0] io_VwirePorts_1_22_0_in,
    input  io_VwirePorts_1_22_0_en,
    output[1:0] io_VwirePorts_1_22_0_out,
    input [1:0] io_VwirePorts_1_21_15_in,
    input  io_VwirePorts_1_21_15_en,
    output[1:0] io_VwirePorts_1_21_15_out,
    input [1:0] io_VwirePorts_1_21_14_in,
    input  io_VwirePorts_1_21_14_en,
    output[1:0] io_VwirePorts_1_21_14_out,
    input [1:0] io_VwirePorts_1_21_13_in,
    input  io_VwirePorts_1_21_13_en,
    output[1:0] io_VwirePorts_1_21_13_out,
    input [1:0] io_VwirePorts_1_21_12_in,
    input  io_VwirePorts_1_21_12_en,
    output[1:0] io_VwirePorts_1_21_12_out,
    input [1:0] io_VwirePorts_1_21_11_in,
    input  io_VwirePorts_1_21_11_en,
    output[1:0] io_VwirePorts_1_21_11_out,
    input [1:0] io_VwirePorts_1_21_10_in,
    input  io_VwirePorts_1_21_10_en,
    output[1:0] io_VwirePorts_1_21_10_out,
    input [1:0] io_VwirePorts_1_21_9_in,
    input  io_VwirePorts_1_21_9_en,
    output[1:0] io_VwirePorts_1_21_9_out,
    input [1:0] io_VwirePorts_1_21_8_in,
    input  io_VwirePorts_1_21_8_en,
    output[1:0] io_VwirePorts_1_21_8_out,
    input [1:0] io_VwirePorts_1_21_7_in,
    input  io_VwirePorts_1_21_7_en,
    output[1:0] io_VwirePorts_1_21_7_out,
    input [1:0] io_VwirePorts_1_21_6_in,
    input  io_VwirePorts_1_21_6_en,
    output[1:0] io_VwirePorts_1_21_6_out,
    input [1:0] io_VwirePorts_1_21_5_in,
    input  io_VwirePorts_1_21_5_en,
    output[1:0] io_VwirePorts_1_21_5_out,
    input [1:0] io_VwirePorts_1_21_4_in,
    input  io_VwirePorts_1_21_4_en,
    output[1:0] io_VwirePorts_1_21_4_out,
    input [1:0] io_VwirePorts_1_21_3_in,
    input  io_VwirePorts_1_21_3_en,
    output[1:0] io_VwirePorts_1_21_3_out,
    input [1:0] io_VwirePorts_1_21_2_in,
    input  io_VwirePorts_1_21_2_en,
    output[1:0] io_VwirePorts_1_21_2_out,
    input [1:0] io_VwirePorts_1_21_1_in,
    input  io_VwirePorts_1_21_1_en,
    output[1:0] io_VwirePorts_1_21_1_out,
    input [1:0] io_VwirePorts_1_21_0_in,
    input  io_VwirePorts_1_21_0_en,
    output[1:0] io_VwirePorts_1_21_0_out,
    input [1:0] io_VwirePorts_1_20_15_in,
    input  io_VwirePorts_1_20_15_en,
    output[1:0] io_VwirePorts_1_20_15_out,
    input [1:0] io_VwirePorts_1_20_14_in,
    input  io_VwirePorts_1_20_14_en,
    output[1:0] io_VwirePorts_1_20_14_out,
    input [1:0] io_VwirePorts_1_20_13_in,
    input  io_VwirePorts_1_20_13_en,
    output[1:0] io_VwirePorts_1_20_13_out,
    input [1:0] io_VwirePorts_1_20_12_in,
    input  io_VwirePorts_1_20_12_en,
    output[1:0] io_VwirePorts_1_20_12_out,
    input [1:0] io_VwirePorts_1_20_11_in,
    input  io_VwirePorts_1_20_11_en,
    output[1:0] io_VwirePorts_1_20_11_out,
    input [1:0] io_VwirePorts_1_20_10_in,
    input  io_VwirePorts_1_20_10_en,
    output[1:0] io_VwirePorts_1_20_10_out,
    input [1:0] io_VwirePorts_1_20_9_in,
    input  io_VwirePorts_1_20_9_en,
    output[1:0] io_VwirePorts_1_20_9_out,
    input [1:0] io_VwirePorts_1_20_8_in,
    input  io_VwirePorts_1_20_8_en,
    output[1:0] io_VwirePorts_1_20_8_out,
    input [1:0] io_VwirePorts_1_20_7_in,
    input  io_VwirePorts_1_20_7_en,
    output[1:0] io_VwirePorts_1_20_7_out,
    input [1:0] io_VwirePorts_1_20_6_in,
    input  io_VwirePorts_1_20_6_en,
    output[1:0] io_VwirePorts_1_20_6_out,
    input [1:0] io_VwirePorts_1_20_5_in,
    input  io_VwirePorts_1_20_5_en,
    output[1:0] io_VwirePorts_1_20_5_out,
    input [1:0] io_VwirePorts_1_20_4_in,
    input  io_VwirePorts_1_20_4_en,
    output[1:0] io_VwirePorts_1_20_4_out,
    input [1:0] io_VwirePorts_1_20_3_in,
    input  io_VwirePorts_1_20_3_en,
    output[1:0] io_VwirePorts_1_20_3_out,
    input [1:0] io_VwirePorts_1_20_2_in,
    input  io_VwirePorts_1_20_2_en,
    output[1:0] io_VwirePorts_1_20_2_out,
    input [1:0] io_VwirePorts_1_20_1_in,
    input  io_VwirePorts_1_20_1_en,
    output[1:0] io_VwirePorts_1_20_1_out,
    input [1:0] io_VwirePorts_1_20_0_in,
    input  io_VwirePorts_1_20_0_en,
    output[1:0] io_VwirePorts_1_20_0_out,
    input [1:0] io_VwirePorts_1_19_15_in,
    input  io_VwirePorts_1_19_15_en,
    output[1:0] io_VwirePorts_1_19_15_out,
    input [1:0] io_VwirePorts_1_19_14_in,
    input  io_VwirePorts_1_19_14_en,
    output[1:0] io_VwirePorts_1_19_14_out,
    input [1:0] io_VwirePorts_1_19_13_in,
    input  io_VwirePorts_1_19_13_en,
    output[1:0] io_VwirePorts_1_19_13_out,
    input [1:0] io_VwirePorts_1_19_12_in,
    input  io_VwirePorts_1_19_12_en,
    output[1:0] io_VwirePorts_1_19_12_out,
    input [1:0] io_VwirePorts_1_19_11_in,
    input  io_VwirePorts_1_19_11_en,
    output[1:0] io_VwirePorts_1_19_11_out,
    input [1:0] io_VwirePorts_1_19_10_in,
    input  io_VwirePorts_1_19_10_en,
    output[1:0] io_VwirePorts_1_19_10_out,
    input [1:0] io_VwirePorts_1_19_9_in,
    input  io_VwirePorts_1_19_9_en,
    output[1:0] io_VwirePorts_1_19_9_out,
    input [1:0] io_VwirePorts_1_19_8_in,
    input  io_VwirePorts_1_19_8_en,
    output[1:0] io_VwirePorts_1_19_8_out,
    input [1:0] io_VwirePorts_1_19_7_in,
    input  io_VwirePorts_1_19_7_en,
    output[1:0] io_VwirePorts_1_19_7_out,
    input [1:0] io_VwirePorts_1_19_6_in,
    input  io_VwirePorts_1_19_6_en,
    output[1:0] io_VwirePorts_1_19_6_out,
    input [1:0] io_VwirePorts_1_19_5_in,
    input  io_VwirePorts_1_19_5_en,
    output[1:0] io_VwirePorts_1_19_5_out,
    input [1:0] io_VwirePorts_1_19_4_in,
    input  io_VwirePorts_1_19_4_en,
    output[1:0] io_VwirePorts_1_19_4_out,
    input [1:0] io_VwirePorts_1_19_3_in,
    input  io_VwirePorts_1_19_3_en,
    output[1:0] io_VwirePorts_1_19_3_out,
    input [1:0] io_VwirePorts_1_19_2_in,
    input  io_VwirePorts_1_19_2_en,
    output[1:0] io_VwirePorts_1_19_2_out,
    input [1:0] io_VwirePorts_1_19_1_in,
    input  io_VwirePorts_1_19_1_en,
    output[1:0] io_VwirePorts_1_19_1_out,
    input [1:0] io_VwirePorts_1_19_0_in,
    input  io_VwirePorts_1_19_0_en,
    output[1:0] io_VwirePorts_1_19_0_out,
    input [1:0] io_VwirePorts_1_18_15_in,
    input  io_VwirePorts_1_18_15_en,
    output[1:0] io_VwirePorts_1_18_15_out,
    input [1:0] io_VwirePorts_1_18_14_in,
    input  io_VwirePorts_1_18_14_en,
    output[1:0] io_VwirePorts_1_18_14_out,
    input [1:0] io_VwirePorts_1_18_13_in,
    input  io_VwirePorts_1_18_13_en,
    output[1:0] io_VwirePorts_1_18_13_out,
    input [1:0] io_VwirePorts_1_18_12_in,
    input  io_VwirePorts_1_18_12_en,
    output[1:0] io_VwirePorts_1_18_12_out,
    input [1:0] io_VwirePorts_1_18_11_in,
    input  io_VwirePorts_1_18_11_en,
    output[1:0] io_VwirePorts_1_18_11_out,
    input [1:0] io_VwirePorts_1_18_10_in,
    input  io_VwirePorts_1_18_10_en,
    output[1:0] io_VwirePorts_1_18_10_out,
    input [1:0] io_VwirePorts_1_18_9_in,
    input  io_VwirePorts_1_18_9_en,
    output[1:0] io_VwirePorts_1_18_9_out,
    input [1:0] io_VwirePorts_1_18_8_in,
    input  io_VwirePorts_1_18_8_en,
    output[1:0] io_VwirePorts_1_18_8_out,
    input [1:0] io_VwirePorts_1_18_7_in,
    input  io_VwirePorts_1_18_7_en,
    output[1:0] io_VwirePorts_1_18_7_out,
    input [1:0] io_VwirePorts_1_18_6_in,
    input  io_VwirePorts_1_18_6_en,
    output[1:0] io_VwirePorts_1_18_6_out,
    input [1:0] io_VwirePorts_1_18_5_in,
    input  io_VwirePorts_1_18_5_en,
    output[1:0] io_VwirePorts_1_18_5_out,
    input [1:0] io_VwirePorts_1_18_4_in,
    input  io_VwirePorts_1_18_4_en,
    output[1:0] io_VwirePorts_1_18_4_out,
    input [1:0] io_VwirePorts_1_18_3_in,
    input  io_VwirePorts_1_18_3_en,
    output[1:0] io_VwirePorts_1_18_3_out,
    input [1:0] io_VwirePorts_1_18_2_in,
    input  io_VwirePorts_1_18_2_en,
    output[1:0] io_VwirePorts_1_18_2_out,
    input [1:0] io_VwirePorts_1_18_1_in,
    input  io_VwirePorts_1_18_1_en,
    output[1:0] io_VwirePorts_1_18_1_out,
    input [1:0] io_VwirePorts_1_18_0_in,
    input  io_VwirePorts_1_18_0_en,
    output[1:0] io_VwirePorts_1_18_0_out,
    input [1:0] io_VwirePorts_1_17_15_in,
    input  io_VwirePorts_1_17_15_en,
    output[1:0] io_VwirePorts_1_17_15_out,
    input [1:0] io_VwirePorts_1_17_14_in,
    input  io_VwirePorts_1_17_14_en,
    output[1:0] io_VwirePorts_1_17_14_out,
    input [1:0] io_VwirePorts_1_17_13_in,
    input  io_VwirePorts_1_17_13_en,
    output[1:0] io_VwirePorts_1_17_13_out,
    input [1:0] io_VwirePorts_1_17_12_in,
    input  io_VwirePorts_1_17_12_en,
    output[1:0] io_VwirePorts_1_17_12_out,
    input [1:0] io_VwirePorts_1_17_11_in,
    input  io_VwirePorts_1_17_11_en,
    output[1:0] io_VwirePorts_1_17_11_out,
    input [1:0] io_VwirePorts_1_17_10_in,
    input  io_VwirePorts_1_17_10_en,
    output[1:0] io_VwirePorts_1_17_10_out,
    input [1:0] io_VwirePorts_1_17_9_in,
    input  io_VwirePorts_1_17_9_en,
    output[1:0] io_VwirePorts_1_17_9_out,
    input [1:0] io_VwirePorts_1_17_8_in,
    input  io_VwirePorts_1_17_8_en,
    output[1:0] io_VwirePorts_1_17_8_out,
    input [1:0] io_VwirePorts_1_17_7_in,
    input  io_VwirePorts_1_17_7_en,
    output[1:0] io_VwirePorts_1_17_7_out,
    input [1:0] io_VwirePorts_1_17_6_in,
    input  io_VwirePorts_1_17_6_en,
    output[1:0] io_VwirePorts_1_17_6_out,
    input [1:0] io_VwirePorts_1_17_5_in,
    input  io_VwirePorts_1_17_5_en,
    output[1:0] io_VwirePorts_1_17_5_out,
    input [1:0] io_VwirePorts_1_17_4_in,
    input  io_VwirePorts_1_17_4_en,
    output[1:0] io_VwirePorts_1_17_4_out,
    input [1:0] io_VwirePorts_1_17_3_in,
    input  io_VwirePorts_1_17_3_en,
    output[1:0] io_VwirePorts_1_17_3_out,
    input [1:0] io_VwirePorts_1_17_2_in,
    input  io_VwirePorts_1_17_2_en,
    output[1:0] io_VwirePorts_1_17_2_out,
    input [1:0] io_VwirePorts_1_17_1_in,
    input  io_VwirePorts_1_17_1_en,
    output[1:0] io_VwirePorts_1_17_1_out,
    input [1:0] io_VwirePorts_1_17_0_in,
    input  io_VwirePorts_1_17_0_en,
    output[1:0] io_VwirePorts_1_17_0_out,
    input [1:0] io_VwirePorts_1_16_15_in,
    input  io_VwirePorts_1_16_15_en,
    output[1:0] io_VwirePorts_1_16_15_out,
    input [1:0] io_VwirePorts_1_16_14_in,
    input  io_VwirePorts_1_16_14_en,
    output[1:0] io_VwirePorts_1_16_14_out,
    input [1:0] io_VwirePorts_1_16_13_in,
    input  io_VwirePorts_1_16_13_en,
    output[1:0] io_VwirePorts_1_16_13_out,
    input [1:0] io_VwirePorts_1_16_12_in,
    input  io_VwirePorts_1_16_12_en,
    output[1:0] io_VwirePorts_1_16_12_out,
    input [1:0] io_VwirePorts_1_16_11_in,
    input  io_VwirePorts_1_16_11_en,
    output[1:0] io_VwirePorts_1_16_11_out,
    input [1:0] io_VwirePorts_1_16_10_in,
    input  io_VwirePorts_1_16_10_en,
    output[1:0] io_VwirePorts_1_16_10_out,
    input [1:0] io_VwirePorts_1_16_9_in,
    input  io_VwirePorts_1_16_9_en,
    output[1:0] io_VwirePorts_1_16_9_out,
    input [1:0] io_VwirePorts_1_16_8_in,
    input  io_VwirePorts_1_16_8_en,
    output[1:0] io_VwirePorts_1_16_8_out,
    input [1:0] io_VwirePorts_1_16_7_in,
    input  io_VwirePorts_1_16_7_en,
    output[1:0] io_VwirePorts_1_16_7_out,
    input [1:0] io_VwirePorts_1_16_6_in,
    input  io_VwirePorts_1_16_6_en,
    output[1:0] io_VwirePorts_1_16_6_out,
    input [1:0] io_VwirePorts_1_16_5_in,
    input  io_VwirePorts_1_16_5_en,
    output[1:0] io_VwirePorts_1_16_5_out,
    input [1:0] io_VwirePorts_1_16_4_in,
    input  io_VwirePorts_1_16_4_en,
    output[1:0] io_VwirePorts_1_16_4_out,
    input [1:0] io_VwirePorts_1_16_3_in,
    input  io_VwirePorts_1_16_3_en,
    output[1:0] io_VwirePorts_1_16_3_out,
    input [1:0] io_VwirePorts_1_16_2_in,
    input  io_VwirePorts_1_16_2_en,
    output[1:0] io_VwirePorts_1_16_2_out,
    input [1:0] io_VwirePorts_1_16_1_in,
    input  io_VwirePorts_1_16_1_en,
    output[1:0] io_VwirePorts_1_16_1_out,
    input [1:0] io_VwirePorts_1_16_0_in,
    input  io_VwirePorts_1_16_0_en,
    output[1:0] io_VwirePorts_1_16_0_out,
    input [1:0] io_VwirePorts_1_15_15_in,
    input  io_VwirePorts_1_15_15_en,
    output[1:0] io_VwirePorts_1_15_15_out,
    input [1:0] io_VwirePorts_1_15_14_in,
    input  io_VwirePorts_1_15_14_en,
    output[1:0] io_VwirePorts_1_15_14_out,
    input [1:0] io_VwirePorts_1_15_13_in,
    input  io_VwirePorts_1_15_13_en,
    output[1:0] io_VwirePorts_1_15_13_out,
    input [1:0] io_VwirePorts_1_15_12_in,
    input  io_VwirePorts_1_15_12_en,
    output[1:0] io_VwirePorts_1_15_12_out,
    input [1:0] io_VwirePorts_1_15_11_in,
    input  io_VwirePorts_1_15_11_en,
    output[1:0] io_VwirePorts_1_15_11_out,
    input [1:0] io_VwirePorts_1_15_10_in,
    input  io_VwirePorts_1_15_10_en,
    output[1:0] io_VwirePorts_1_15_10_out,
    input [1:0] io_VwirePorts_1_15_9_in,
    input  io_VwirePorts_1_15_9_en,
    output[1:0] io_VwirePorts_1_15_9_out,
    input [1:0] io_VwirePorts_1_15_8_in,
    input  io_VwirePorts_1_15_8_en,
    output[1:0] io_VwirePorts_1_15_8_out,
    input [1:0] io_VwirePorts_1_15_7_in,
    input  io_VwirePorts_1_15_7_en,
    output[1:0] io_VwirePorts_1_15_7_out,
    input [1:0] io_VwirePorts_1_15_6_in,
    input  io_VwirePorts_1_15_6_en,
    output[1:0] io_VwirePorts_1_15_6_out,
    input [1:0] io_VwirePorts_1_15_5_in,
    input  io_VwirePorts_1_15_5_en,
    output[1:0] io_VwirePorts_1_15_5_out,
    input [1:0] io_VwirePorts_1_15_4_in,
    input  io_VwirePorts_1_15_4_en,
    output[1:0] io_VwirePorts_1_15_4_out,
    input [1:0] io_VwirePorts_1_15_3_in,
    input  io_VwirePorts_1_15_3_en,
    output[1:0] io_VwirePorts_1_15_3_out,
    input [1:0] io_VwirePorts_1_15_2_in,
    input  io_VwirePorts_1_15_2_en,
    output[1:0] io_VwirePorts_1_15_2_out,
    input [1:0] io_VwirePorts_1_15_1_in,
    input  io_VwirePorts_1_15_1_en,
    output[1:0] io_VwirePorts_1_15_1_out,
    input [1:0] io_VwirePorts_1_15_0_in,
    input  io_VwirePorts_1_15_0_en,
    output[1:0] io_VwirePorts_1_15_0_out,
    input [1:0] io_VwirePorts_1_14_15_in,
    input  io_VwirePorts_1_14_15_en,
    output[1:0] io_VwirePorts_1_14_15_out,
    input [1:0] io_VwirePorts_1_14_14_in,
    input  io_VwirePorts_1_14_14_en,
    output[1:0] io_VwirePorts_1_14_14_out,
    input [1:0] io_VwirePorts_1_14_13_in,
    input  io_VwirePorts_1_14_13_en,
    output[1:0] io_VwirePorts_1_14_13_out,
    input [1:0] io_VwirePorts_1_14_12_in,
    input  io_VwirePorts_1_14_12_en,
    output[1:0] io_VwirePorts_1_14_12_out,
    input [1:0] io_VwirePorts_1_14_11_in,
    input  io_VwirePorts_1_14_11_en,
    output[1:0] io_VwirePorts_1_14_11_out,
    input [1:0] io_VwirePorts_1_14_10_in,
    input  io_VwirePorts_1_14_10_en,
    output[1:0] io_VwirePorts_1_14_10_out,
    input [1:0] io_VwirePorts_1_14_9_in,
    input  io_VwirePorts_1_14_9_en,
    output[1:0] io_VwirePorts_1_14_9_out,
    input [1:0] io_VwirePorts_1_14_8_in,
    input  io_VwirePorts_1_14_8_en,
    output[1:0] io_VwirePorts_1_14_8_out,
    input [1:0] io_VwirePorts_1_14_7_in,
    input  io_VwirePorts_1_14_7_en,
    output[1:0] io_VwirePorts_1_14_7_out,
    input [1:0] io_VwirePorts_1_14_6_in,
    input  io_VwirePorts_1_14_6_en,
    output[1:0] io_VwirePorts_1_14_6_out,
    input [1:0] io_VwirePorts_1_14_5_in,
    input  io_VwirePorts_1_14_5_en,
    output[1:0] io_VwirePorts_1_14_5_out,
    input [1:0] io_VwirePorts_1_14_4_in,
    input  io_VwirePorts_1_14_4_en,
    output[1:0] io_VwirePorts_1_14_4_out,
    input [1:0] io_VwirePorts_1_14_3_in,
    input  io_VwirePorts_1_14_3_en,
    output[1:0] io_VwirePorts_1_14_3_out,
    input [1:0] io_VwirePorts_1_14_2_in,
    input  io_VwirePorts_1_14_2_en,
    output[1:0] io_VwirePorts_1_14_2_out,
    input [1:0] io_VwirePorts_1_14_1_in,
    input  io_VwirePorts_1_14_1_en,
    output[1:0] io_VwirePorts_1_14_1_out,
    input [1:0] io_VwirePorts_1_14_0_in,
    input  io_VwirePorts_1_14_0_en,
    output[1:0] io_VwirePorts_1_14_0_out,
    input [1:0] io_VwirePorts_1_13_15_in,
    input  io_VwirePorts_1_13_15_en,
    output[1:0] io_VwirePorts_1_13_15_out,
    input [1:0] io_VwirePorts_1_13_14_in,
    input  io_VwirePorts_1_13_14_en,
    output[1:0] io_VwirePorts_1_13_14_out,
    input [1:0] io_VwirePorts_1_13_13_in,
    input  io_VwirePorts_1_13_13_en,
    output[1:0] io_VwirePorts_1_13_13_out,
    input [1:0] io_VwirePorts_1_13_12_in,
    input  io_VwirePorts_1_13_12_en,
    output[1:0] io_VwirePorts_1_13_12_out,
    input [1:0] io_VwirePorts_1_13_11_in,
    input  io_VwirePorts_1_13_11_en,
    output[1:0] io_VwirePorts_1_13_11_out,
    input [1:0] io_VwirePorts_1_13_10_in,
    input  io_VwirePorts_1_13_10_en,
    output[1:0] io_VwirePorts_1_13_10_out,
    input [1:0] io_VwirePorts_1_13_9_in,
    input  io_VwirePorts_1_13_9_en,
    output[1:0] io_VwirePorts_1_13_9_out,
    input [1:0] io_VwirePorts_1_13_8_in,
    input  io_VwirePorts_1_13_8_en,
    output[1:0] io_VwirePorts_1_13_8_out,
    input [1:0] io_VwirePorts_1_13_7_in,
    input  io_VwirePorts_1_13_7_en,
    output[1:0] io_VwirePorts_1_13_7_out,
    input [1:0] io_VwirePorts_1_13_6_in,
    input  io_VwirePorts_1_13_6_en,
    output[1:0] io_VwirePorts_1_13_6_out,
    input [1:0] io_VwirePorts_1_13_5_in,
    input  io_VwirePorts_1_13_5_en,
    output[1:0] io_VwirePorts_1_13_5_out,
    input [1:0] io_VwirePorts_1_13_4_in,
    input  io_VwirePorts_1_13_4_en,
    output[1:0] io_VwirePorts_1_13_4_out,
    input [1:0] io_VwirePorts_1_13_3_in,
    input  io_VwirePorts_1_13_3_en,
    output[1:0] io_VwirePorts_1_13_3_out,
    input [1:0] io_VwirePorts_1_13_2_in,
    input  io_VwirePorts_1_13_2_en,
    output[1:0] io_VwirePorts_1_13_2_out,
    input [1:0] io_VwirePorts_1_13_1_in,
    input  io_VwirePorts_1_13_1_en,
    output[1:0] io_VwirePorts_1_13_1_out,
    input [1:0] io_VwirePorts_1_13_0_in,
    input  io_VwirePorts_1_13_0_en,
    output[1:0] io_VwirePorts_1_13_0_out,
    input [1:0] io_VwirePorts_1_12_15_in,
    input  io_VwirePorts_1_12_15_en,
    output[1:0] io_VwirePorts_1_12_15_out,
    input [1:0] io_VwirePorts_1_12_14_in,
    input  io_VwirePorts_1_12_14_en,
    output[1:0] io_VwirePorts_1_12_14_out,
    input [1:0] io_VwirePorts_1_12_13_in,
    input  io_VwirePorts_1_12_13_en,
    output[1:0] io_VwirePorts_1_12_13_out,
    input [1:0] io_VwirePorts_1_12_12_in,
    input  io_VwirePorts_1_12_12_en,
    output[1:0] io_VwirePorts_1_12_12_out,
    input [1:0] io_VwirePorts_1_12_11_in,
    input  io_VwirePorts_1_12_11_en,
    output[1:0] io_VwirePorts_1_12_11_out,
    input [1:0] io_VwirePorts_1_12_10_in,
    input  io_VwirePorts_1_12_10_en,
    output[1:0] io_VwirePorts_1_12_10_out,
    input [1:0] io_VwirePorts_1_12_9_in,
    input  io_VwirePorts_1_12_9_en,
    output[1:0] io_VwirePorts_1_12_9_out,
    input [1:0] io_VwirePorts_1_12_8_in,
    input  io_VwirePorts_1_12_8_en,
    output[1:0] io_VwirePorts_1_12_8_out,
    input [1:0] io_VwirePorts_1_12_7_in,
    input  io_VwirePorts_1_12_7_en,
    output[1:0] io_VwirePorts_1_12_7_out,
    input [1:0] io_VwirePorts_1_12_6_in,
    input  io_VwirePorts_1_12_6_en,
    output[1:0] io_VwirePorts_1_12_6_out,
    input [1:0] io_VwirePorts_1_12_5_in,
    input  io_VwirePorts_1_12_5_en,
    output[1:0] io_VwirePorts_1_12_5_out,
    input [1:0] io_VwirePorts_1_12_4_in,
    input  io_VwirePorts_1_12_4_en,
    output[1:0] io_VwirePorts_1_12_4_out,
    input [1:0] io_VwirePorts_1_12_3_in,
    input  io_VwirePorts_1_12_3_en,
    output[1:0] io_VwirePorts_1_12_3_out,
    input [1:0] io_VwirePorts_1_12_2_in,
    input  io_VwirePorts_1_12_2_en,
    output[1:0] io_VwirePorts_1_12_2_out,
    input [1:0] io_VwirePorts_1_12_1_in,
    input  io_VwirePorts_1_12_1_en,
    output[1:0] io_VwirePorts_1_12_1_out,
    input [1:0] io_VwirePorts_1_12_0_in,
    input  io_VwirePorts_1_12_0_en,
    output[1:0] io_VwirePorts_1_12_0_out,
    input [1:0] io_VwirePorts_1_11_15_in,
    input  io_VwirePorts_1_11_15_en,
    output[1:0] io_VwirePorts_1_11_15_out,
    input [1:0] io_VwirePorts_1_11_14_in,
    input  io_VwirePorts_1_11_14_en,
    output[1:0] io_VwirePorts_1_11_14_out,
    input [1:0] io_VwirePorts_1_11_13_in,
    input  io_VwirePorts_1_11_13_en,
    output[1:0] io_VwirePorts_1_11_13_out,
    input [1:0] io_VwirePorts_1_11_12_in,
    input  io_VwirePorts_1_11_12_en,
    output[1:0] io_VwirePorts_1_11_12_out,
    input [1:0] io_VwirePorts_1_11_11_in,
    input  io_VwirePorts_1_11_11_en,
    output[1:0] io_VwirePorts_1_11_11_out,
    input [1:0] io_VwirePorts_1_11_10_in,
    input  io_VwirePorts_1_11_10_en,
    output[1:0] io_VwirePorts_1_11_10_out,
    input [1:0] io_VwirePorts_1_11_9_in,
    input  io_VwirePorts_1_11_9_en,
    output[1:0] io_VwirePorts_1_11_9_out,
    input [1:0] io_VwirePorts_1_11_8_in,
    input  io_VwirePorts_1_11_8_en,
    output[1:0] io_VwirePorts_1_11_8_out,
    input [1:0] io_VwirePorts_1_11_7_in,
    input  io_VwirePorts_1_11_7_en,
    output[1:0] io_VwirePorts_1_11_7_out,
    input [1:0] io_VwirePorts_1_11_6_in,
    input  io_VwirePorts_1_11_6_en,
    output[1:0] io_VwirePorts_1_11_6_out,
    input [1:0] io_VwirePorts_1_11_5_in,
    input  io_VwirePorts_1_11_5_en,
    output[1:0] io_VwirePorts_1_11_5_out,
    input [1:0] io_VwirePorts_1_11_4_in,
    input  io_VwirePorts_1_11_4_en,
    output[1:0] io_VwirePorts_1_11_4_out,
    input [1:0] io_VwirePorts_1_11_3_in,
    input  io_VwirePorts_1_11_3_en,
    output[1:0] io_VwirePorts_1_11_3_out,
    input [1:0] io_VwirePorts_1_11_2_in,
    input  io_VwirePorts_1_11_2_en,
    output[1:0] io_VwirePorts_1_11_2_out,
    input [1:0] io_VwirePorts_1_11_1_in,
    input  io_VwirePorts_1_11_1_en,
    output[1:0] io_VwirePorts_1_11_1_out,
    input [1:0] io_VwirePorts_1_11_0_in,
    input  io_VwirePorts_1_11_0_en,
    output[1:0] io_VwirePorts_1_11_0_out,
    input [1:0] io_VwirePorts_1_10_15_in,
    input  io_VwirePorts_1_10_15_en,
    output[1:0] io_VwirePorts_1_10_15_out,
    input [1:0] io_VwirePorts_1_10_14_in,
    input  io_VwirePorts_1_10_14_en,
    output[1:0] io_VwirePorts_1_10_14_out,
    input [1:0] io_VwirePorts_1_10_13_in,
    input  io_VwirePorts_1_10_13_en,
    output[1:0] io_VwirePorts_1_10_13_out,
    input [1:0] io_VwirePorts_1_10_12_in,
    input  io_VwirePorts_1_10_12_en,
    output[1:0] io_VwirePorts_1_10_12_out,
    input [1:0] io_VwirePorts_1_10_11_in,
    input  io_VwirePorts_1_10_11_en,
    output[1:0] io_VwirePorts_1_10_11_out,
    input [1:0] io_VwirePorts_1_10_10_in,
    input  io_VwirePorts_1_10_10_en,
    output[1:0] io_VwirePorts_1_10_10_out,
    input [1:0] io_VwirePorts_1_10_9_in,
    input  io_VwirePorts_1_10_9_en,
    output[1:0] io_VwirePorts_1_10_9_out,
    input [1:0] io_VwirePorts_1_10_8_in,
    input  io_VwirePorts_1_10_8_en,
    output[1:0] io_VwirePorts_1_10_8_out,
    input [1:0] io_VwirePorts_1_10_7_in,
    input  io_VwirePorts_1_10_7_en,
    output[1:0] io_VwirePorts_1_10_7_out,
    input [1:0] io_VwirePorts_1_10_6_in,
    input  io_VwirePorts_1_10_6_en,
    output[1:0] io_VwirePorts_1_10_6_out,
    input [1:0] io_VwirePorts_1_10_5_in,
    input  io_VwirePorts_1_10_5_en,
    output[1:0] io_VwirePorts_1_10_5_out,
    input [1:0] io_VwirePorts_1_10_4_in,
    input  io_VwirePorts_1_10_4_en,
    output[1:0] io_VwirePorts_1_10_4_out,
    input [1:0] io_VwirePorts_1_10_3_in,
    input  io_VwirePorts_1_10_3_en,
    output[1:0] io_VwirePorts_1_10_3_out,
    input [1:0] io_VwirePorts_1_10_2_in,
    input  io_VwirePorts_1_10_2_en,
    output[1:0] io_VwirePorts_1_10_2_out,
    input [1:0] io_VwirePorts_1_10_1_in,
    input  io_VwirePorts_1_10_1_en,
    output[1:0] io_VwirePorts_1_10_1_out,
    input [1:0] io_VwirePorts_1_10_0_in,
    input  io_VwirePorts_1_10_0_en,
    output[1:0] io_VwirePorts_1_10_0_out,
    input [1:0] io_VwirePorts_1_9_15_in,
    input  io_VwirePorts_1_9_15_en,
    output[1:0] io_VwirePorts_1_9_15_out,
    input [1:0] io_VwirePorts_1_9_14_in,
    input  io_VwirePorts_1_9_14_en,
    output[1:0] io_VwirePorts_1_9_14_out,
    input [1:0] io_VwirePorts_1_9_13_in,
    input  io_VwirePorts_1_9_13_en,
    output[1:0] io_VwirePorts_1_9_13_out,
    input [1:0] io_VwirePorts_1_9_12_in,
    input  io_VwirePorts_1_9_12_en,
    output[1:0] io_VwirePorts_1_9_12_out,
    input [1:0] io_VwirePorts_1_9_11_in,
    input  io_VwirePorts_1_9_11_en,
    output[1:0] io_VwirePorts_1_9_11_out,
    input [1:0] io_VwirePorts_1_9_10_in,
    input  io_VwirePorts_1_9_10_en,
    output[1:0] io_VwirePorts_1_9_10_out,
    input [1:0] io_VwirePorts_1_9_9_in,
    input  io_VwirePorts_1_9_9_en,
    output[1:0] io_VwirePorts_1_9_9_out,
    input [1:0] io_VwirePorts_1_9_8_in,
    input  io_VwirePorts_1_9_8_en,
    output[1:0] io_VwirePorts_1_9_8_out,
    input [1:0] io_VwirePorts_1_9_7_in,
    input  io_VwirePorts_1_9_7_en,
    output[1:0] io_VwirePorts_1_9_7_out,
    input [1:0] io_VwirePorts_1_9_6_in,
    input  io_VwirePorts_1_9_6_en,
    output[1:0] io_VwirePorts_1_9_6_out,
    input [1:0] io_VwirePorts_1_9_5_in,
    input  io_VwirePorts_1_9_5_en,
    output[1:0] io_VwirePorts_1_9_5_out,
    input [1:0] io_VwirePorts_1_9_4_in,
    input  io_VwirePorts_1_9_4_en,
    output[1:0] io_VwirePorts_1_9_4_out,
    input [1:0] io_VwirePorts_1_9_3_in,
    input  io_VwirePorts_1_9_3_en,
    output[1:0] io_VwirePorts_1_9_3_out,
    input [1:0] io_VwirePorts_1_9_2_in,
    input  io_VwirePorts_1_9_2_en,
    output[1:0] io_VwirePorts_1_9_2_out,
    input [1:0] io_VwirePorts_1_9_1_in,
    input  io_VwirePorts_1_9_1_en,
    output[1:0] io_VwirePorts_1_9_1_out,
    input [1:0] io_VwirePorts_1_9_0_in,
    input  io_VwirePorts_1_9_0_en,
    output[1:0] io_VwirePorts_1_9_0_out,
    input [1:0] io_VwirePorts_1_8_15_in,
    input  io_VwirePorts_1_8_15_en,
    output[1:0] io_VwirePorts_1_8_15_out,
    input [1:0] io_VwirePorts_1_8_14_in,
    input  io_VwirePorts_1_8_14_en,
    output[1:0] io_VwirePorts_1_8_14_out,
    input [1:0] io_VwirePorts_1_8_13_in,
    input  io_VwirePorts_1_8_13_en,
    output[1:0] io_VwirePorts_1_8_13_out,
    input [1:0] io_VwirePorts_1_8_12_in,
    input  io_VwirePorts_1_8_12_en,
    output[1:0] io_VwirePorts_1_8_12_out,
    input [1:0] io_VwirePorts_1_8_11_in,
    input  io_VwirePorts_1_8_11_en,
    output[1:0] io_VwirePorts_1_8_11_out,
    input [1:0] io_VwirePorts_1_8_10_in,
    input  io_VwirePorts_1_8_10_en,
    output[1:0] io_VwirePorts_1_8_10_out,
    input [1:0] io_VwirePorts_1_8_9_in,
    input  io_VwirePorts_1_8_9_en,
    output[1:0] io_VwirePorts_1_8_9_out,
    input [1:0] io_VwirePorts_1_8_8_in,
    input  io_VwirePorts_1_8_8_en,
    output[1:0] io_VwirePorts_1_8_8_out,
    input [1:0] io_VwirePorts_1_8_7_in,
    input  io_VwirePorts_1_8_7_en,
    output[1:0] io_VwirePorts_1_8_7_out,
    input [1:0] io_VwirePorts_1_8_6_in,
    input  io_VwirePorts_1_8_6_en,
    output[1:0] io_VwirePorts_1_8_6_out,
    input [1:0] io_VwirePorts_1_8_5_in,
    input  io_VwirePorts_1_8_5_en,
    output[1:0] io_VwirePorts_1_8_5_out,
    input [1:0] io_VwirePorts_1_8_4_in,
    input  io_VwirePorts_1_8_4_en,
    output[1:0] io_VwirePorts_1_8_4_out,
    input [1:0] io_VwirePorts_1_8_3_in,
    input  io_VwirePorts_1_8_3_en,
    output[1:0] io_VwirePorts_1_8_3_out,
    input [1:0] io_VwirePorts_1_8_2_in,
    input  io_VwirePorts_1_8_2_en,
    output[1:0] io_VwirePorts_1_8_2_out,
    input [1:0] io_VwirePorts_1_8_1_in,
    input  io_VwirePorts_1_8_1_en,
    output[1:0] io_VwirePorts_1_8_1_out,
    input [1:0] io_VwirePorts_1_8_0_in,
    input  io_VwirePorts_1_8_0_en,
    output[1:0] io_VwirePorts_1_8_0_out,
    input [1:0] io_VwirePorts_1_7_15_in,
    input  io_VwirePorts_1_7_15_en,
    output[1:0] io_VwirePorts_1_7_15_out,
    input [1:0] io_VwirePorts_1_7_14_in,
    input  io_VwirePorts_1_7_14_en,
    output[1:0] io_VwirePorts_1_7_14_out,
    input [1:0] io_VwirePorts_1_7_13_in,
    input  io_VwirePorts_1_7_13_en,
    output[1:0] io_VwirePorts_1_7_13_out,
    input [1:0] io_VwirePorts_1_7_12_in,
    input  io_VwirePorts_1_7_12_en,
    output[1:0] io_VwirePorts_1_7_12_out,
    input [1:0] io_VwirePorts_1_7_11_in,
    input  io_VwirePorts_1_7_11_en,
    output[1:0] io_VwirePorts_1_7_11_out,
    input [1:0] io_VwirePorts_1_7_10_in,
    input  io_VwirePorts_1_7_10_en,
    output[1:0] io_VwirePorts_1_7_10_out,
    input [1:0] io_VwirePorts_1_7_9_in,
    input  io_VwirePorts_1_7_9_en,
    output[1:0] io_VwirePorts_1_7_9_out,
    input [1:0] io_VwirePorts_1_7_8_in,
    input  io_VwirePorts_1_7_8_en,
    output[1:0] io_VwirePorts_1_7_8_out,
    input [1:0] io_VwirePorts_1_7_7_in,
    input  io_VwirePorts_1_7_7_en,
    output[1:0] io_VwirePorts_1_7_7_out,
    input [1:0] io_VwirePorts_1_7_6_in,
    input  io_VwirePorts_1_7_6_en,
    output[1:0] io_VwirePorts_1_7_6_out,
    input [1:0] io_VwirePorts_1_7_5_in,
    input  io_VwirePorts_1_7_5_en,
    output[1:0] io_VwirePorts_1_7_5_out,
    input [1:0] io_VwirePorts_1_7_4_in,
    input  io_VwirePorts_1_7_4_en,
    output[1:0] io_VwirePorts_1_7_4_out,
    input [1:0] io_VwirePorts_1_7_3_in,
    input  io_VwirePorts_1_7_3_en,
    output[1:0] io_VwirePorts_1_7_3_out,
    input [1:0] io_VwirePorts_1_7_2_in,
    input  io_VwirePorts_1_7_2_en,
    output[1:0] io_VwirePorts_1_7_2_out,
    input [1:0] io_VwirePorts_1_7_1_in,
    input  io_VwirePorts_1_7_1_en,
    output[1:0] io_VwirePorts_1_7_1_out,
    input [1:0] io_VwirePorts_1_7_0_in,
    input  io_VwirePorts_1_7_0_en,
    output[1:0] io_VwirePorts_1_7_0_out,
    input [1:0] io_VwirePorts_1_6_15_in,
    input  io_VwirePorts_1_6_15_en,
    output[1:0] io_VwirePorts_1_6_15_out,
    input [1:0] io_VwirePorts_1_6_14_in,
    input  io_VwirePorts_1_6_14_en,
    output[1:0] io_VwirePorts_1_6_14_out,
    input [1:0] io_VwirePorts_1_6_13_in,
    input  io_VwirePorts_1_6_13_en,
    output[1:0] io_VwirePorts_1_6_13_out,
    input [1:0] io_VwirePorts_1_6_12_in,
    input  io_VwirePorts_1_6_12_en,
    output[1:0] io_VwirePorts_1_6_12_out,
    input [1:0] io_VwirePorts_1_6_11_in,
    input  io_VwirePorts_1_6_11_en,
    output[1:0] io_VwirePorts_1_6_11_out,
    input [1:0] io_VwirePorts_1_6_10_in,
    input  io_VwirePorts_1_6_10_en,
    output[1:0] io_VwirePorts_1_6_10_out,
    input [1:0] io_VwirePorts_1_6_9_in,
    input  io_VwirePorts_1_6_9_en,
    output[1:0] io_VwirePorts_1_6_9_out,
    input [1:0] io_VwirePorts_1_6_8_in,
    input  io_VwirePorts_1_6_8_en,
    output[1:0] io_VwirePorts_1_6_8_out,
    input [1:0] io_VwirePorts_1_6_7_in,
    input  io_VwirePorts_1_6_7_en,
    output[1:0] io_VwirePorts_1_6_7_out,
    input [1:0] io_VwirePorts_1_6_6_in,
    input  io_VwirePorts_1_6_6_en,
    output[1:0] io_VwirePorts_1_6_6_out,
    input [1:0] io_VwirePorts_1_6_5_in,
    input  io_VwirePorts_1_6_5_en,
    output[1:0] io_VwirePorts_1_6_5_out,
    input [1:0] io_VwirePorts_1_6_4_in,
    input  io_VwirePorts_1_6_4_en,
    output[1:0] io_VwirePorts_1_6_4_out,
    input [1:0] io_VwirePorts_1_6_3_in,
    input  io_VwirePorts_1_6_3_en,
    output[1:0] io_VwirePorts_1_6_3_out,
    input [1:0] io_VwirePorts_1_6_2_in,
    input  io_VwirePorts_1_6_2_en,
    output[1:0] io_VwirePorts_1_6_2_out,
    input [1:0] io_VwirePorts_1_6_1_in,
    input  io_VwirePorts_1_6_1_en,
    output[1:0] io_VwirePorts_1_6_1_out,
    input [1:0] io_VwirePorts_1_6_0_in,
    input  io_VwirePorts_1_6_0_en,
    output[1:0] io_VwirePorts_1_6_0_out,
    input [1:0] io_VwirePorts_1_5_15_in,
    input  io_VwirePorts_1_5_15_en,
    output[1:0] io_VwirePorts_1_5_15_out,
    input [1:0] io_VwirePorts_1_5_14_in,
    input  io_VwirePorts_1_5_14_en,
    output[1:0] io_VwirePorts_1_5_14_out,
    input [1:0] io_VwirePorts_1_5_13_in,
    input  io_VwirePorts_1_5_13_en,
    output[1:0] io_VwirePorts_1_5_13_out,
    input [1:0] io_VwirePorts_1_5_12_in,
    input  io_VwirePorts_1_5_12_en,
    output[1:0] io_VwirePorts_1_5_12_out,
    input [1:0] io_VwirePorts_1_5_11_in,
    input  io_VwirePorts_1_5_11_en,
    output[1:0] io_VwirePorts_1_5_11_out,
    input [1:0] io_VwirePorts_1_5_10_in,
    input  io_VwirePorts_1_5_10_en,
    output[1:0] io_VwirePorts_1_5_10_out,
    input [1:0] io_VwirePorts_1_5_9_in,
    input  io_VwirePorts_1_5_9_en,
    output[1:0] io_VwirePorts_1_5_9_out,
    input [1:0] io_VwirePorts_1_5_8_in,
    input  io_VwirePorts_1_5_8_en,
    output[1:0] io_VwirePorts_1_5_8_out,
    input [1:0] io_VwirePorts_1_5_7_in,
    input  io_VwirePorts_1_5_7_en,
    output[1:0] io_VwirePorts_1_5_7_out,
    input [1:0] io_VwirePorts_1_5_6_in,
    input  io_VwirePorts_1_5_6_en,
    output[1:0] io_VwirePorts_1_5_6_out,
    input [1:0] io_VwirePorts_1_5_5_in,
    input  io_VwirePorts_1_5_5_en,
    output[1:0] io_VwirePorts_1_5_5_out,
    input [1:0] io_VwirePorts_1_5_4_in,
    input  io_VwirePorts_1_5_4_en,
    output[1:0] io_VwirePorts_1_5_4_out,
    input [1:0] io_VwirePorts_1_5_3_in,
    input  io_VwirePorts_1_5_3_en,
    output[1:0] io_VwirePorts_1_5_3_out,
    input [1:0] io_VwirePorts_1_5_2_in,
    input  io_VwirePorts_1_5_2_en,
    output[1:0] io_VwirePorts_1_5_2_out,
    input [1:0] io_VwirePorts_1_5_1_in,
    input  io_VwirePorts_1_5_1_en,
    output[1:0] io_VwirePorts_1_5_1_out,
    input [1:0] io_VwirePorts_1_5_0_in,
    input  io_VwirePorts_1_5_0_en,
    output[1:0] io_VwirePorts_1_5_0_out,
    input [1:0] io_VwirePorts_1_4_15_in,
    input  io_VwirePorts_1_4_15_en,
    output[1:0] io_VwirePorts_1_4_15_out,
    input [1:0] io_VwirePorts_1_4_14_in,
    input  io_VwirePorts_1_4_14_en,
    output[1:0] io_VwirePorts_1_4_14_out,
    input [1:0] io_VwirePorts_1_4_13_in,
    input  io_VwirePorts_1_4_13_en,
    output[1:0] io_VwirePorts_1_4_13_out,
    input [1:0] io_VwirePorts_1_4_12_in,
    input  io_VwirePorts_1_4_12_en,
    output[1:0] io_VwirePorts_1_4_12_out,
    input [1:0] io_VwirePorts_1_4_11_in,
    input  io_VwirePorts_1_4_11_en,
    output[1:0] io_VwirePorts_1_4_11_out,
    input [1:0] io_VwirePorts_1_4_10_in,
    input  io_VwirePorts_1_4_10_en,
    output[1:0] io_VwirePorts_1_4_10_out,
    input [1:0] io_VwirePorts_1_4_9_in,
    input  io_VwirePorts_1_4_9_en,
    output[1:0] io_VwirePorts_1_4_9_out,
    input [1:0] io_VwirePorts_1_4_8_in,
    input  io_VwirePorts_1_4_8_en,
    output[1:0] io_VwirePorts_1_4_8_out,
    input [1:0] io_VwirePorts_1_4_7_in,
    input  io_VwirePorts_1_4_7_en,
    output[1:0] io_VwirePorts_1_4_7_out,
    input [1:0] io_VwirePorts_1_4_6_in,
    input  io_VwirePorts_1_4_6_en,
    output[1:0] io_VwirePorts_1_4_6_out,
    input [1:0] io_VwirePorts_1_4_5_in,
    input  io_VwirePorts_1_4_5_en,
    output[1:0] io_VwirePorts_1_4_5_out,
    input [1:0] io_VwirePorts_1_4_4_in,
    input  io_VwirePorts_1_4_4_en,
    output[1:0] io_VwirePorts_1_4_4_out,
    input [1:0] io_VwirePorts_1_4_3_in,
    input  io_VwirePorts_1_4_3_en,
    output[1:0] io_VwirePorts_1_4_3_out,
    input [1:0] io_VwirePorts_1_4_2_in,
    input  io_VwirePorts_1_4_2_en,
    output[1:0] io_VwirePorts_1_4_2_out,
    input [1:0] io_VwirePorts_1_4_1_in,
    input  io_VwirePorts_1_4_1_en,
    output[1:0] io_VwirePorts_1_4_1_out,
    input [1:0] io_VwirePorts_1_4_0_in,
    input  io_VwirePorts_1_4_0_en,
    output[1:0] io_VwirePorts_1_4_0_out,
    input [1:0] io_VwirePorts_1_3_15_in,
    input  io_VwirePorts_1_3_15_en,
    output[1:0] io_VwirePorts_1_3_15_out,
    input [1:0] io_VwirePorts_1_3_14_in,
    input  io_VwirePorts_1_3_14_en,
    output[1:0] io_VwirePorts_1_3_14_out,
    input [1:0] io_VwirePorts_1_3_13_in,
    input  io_VwirePorts_1_3_13_en,
    output[1:0] io_VwirePorts_1_3_13_out,
    input [1:0] io_VwirePorts_1_3_12_in,
    input  io_VwirePorts_1_3_12_en,
    output[1:0] io_VwirePorts_1_3_12_out,
    input [1:0] io_VwirePorts_1_3_11_in,
    input  io_VwirePorts_1_3_11_en,
    output[1:0] io_VwirePorts_1_3_11_out,
    input [1:0] io_VwirePorts_1_3_10_in,
    input  io_VwirePorts_1_3_10_en,
    output[1:0] io_VwirePorts_1_3_10_out,
    input [1:0] io_VwirePorts_1_3_9_in,
    input  io_VwirePorts_1_3_9_en,
    output[1:0] io_VwirePorts_1_3_9_out,
    input [1:0] io_VwirePorts_1_3_8_in,
    input  io_VwirePorts_1_3_8_en,
    output[1:0] io_VwirePorts_1_3_8_out,
    input [1:0] io_VwirePorts_1_3_7_in,
    input  io_VwirePorts_1_3_7_en,
    output[1:0] io_VwirePorts_1_3_7_out,
    input [1:0] io_VwirePorts_1_3_6_in,
    input  io_VwirePorts_1_3_6_en,
    output[1:0] io_VwirePorts_1_3_6_out,
    input [1:0] io_VwirePorts_1_3_5_in,
    input  io_VwirePorts_1_3_5_en,
    output[1:0] io_VwirePorts_1_3_5_out,
    input [1:0] io_VwirePorts_1_3_4_in,
    input  io_VwirePorts_1_3_4_en,
    output[1:0] io_VwirePorts_1_3_4_out,
    input [1:0] io_VwirePorts_1_3_3_in,
    input  io_VwirePorts_1_3_3_en,
    output[1:0] io_VwirePorts_1_3_3_out,
    input [1:0] io_VwirePorts_1_3_2_in,
    input  io_VwirePorts_1_3_2_en,
    output[1:0] io_VwirePorts_1_3_2_out,
    input [1:0] io_VwirePorts_1_3_1_in,
    input  io_VwirePorts_1_3_1_en,
    output[1:0] io_VwirePorts_1_3_1_out,
    input [1:0] io_VwirePorts_1_3_0_in,
    input  io_VwirePorts_1_3_0_en,
    output[1:0] io_VwirePorts_1_3_0_out,
    input [1:0] io_VwirePorts_1_2_15_in,
    input  io_VwirePorts_1_2_15_en,
    output[1:0] io_VwirePorts_1_2_15_out,
    input [1:0] io_VwirePorts_1_2_14_in,
    input  io_VwirePorts_1_2_14_en,
    output[1:0] io_VwirePorts_1_2_14_out,
    input [1:0] io_VwirePorts_1_2_13_in,
    input  io_VwirePorts_1_2_13_en,
    output[1:0] io_VwirePorts_1_2_13_out,
    input [1:0] io_VwirePorts_1_2_12_in,
    input  io_VwirePorts_1_2_12_en,
    output[1:0] io_VwirePorts_1_2_12_out,
    input [1:0] io_VwirePorts_1_2_11_in,
    input  io_VwirePorts_1_2_11_en,
    output[1:0] io_VwirePorts_1_2_11_out,
    input [1:0] io_VwirePorts_1_2_10_in,
    input  io_VwirePorts_1_2_10_en,
    output[1:0] io_VwirePorts_1_2_10_out,
    input [1:0] io_VwirePorts_1_2_9_in,
    input  io_VwirePorts_1_2_9_en,
    output[1:0] io_VwirePorts_1_2_9_out,
    input [1:0] io_VwirePorts_1_2_8_in,
    input  io_VwirePorts_1_2_8_en,
    output[1:0] io_VwirePorts_1_2_8_out,
    input [1:0] io_VwirePorts_1_2_7_in,
    input  io_VwirePorts_1_2_7_en,
    output[1:0] io_VwirePorts_1_2_7_out,
    input [1:0] io_VwirePorts_1_2_6_in,
    input  io_VwirePorts_1_2_6_en,
    output[1:0] io_VwirePorts_1_2_6_out,
    input [1:0] io_VwirePorts_1_2_5_in,
    input  io_VwirePorts_1_2_5_en,
    output[1:0] io_VwirePorts_1_2_5_out,
    input [1:0] io_VwirePorts_1_2_4_in,
    input  io_VwirePorts_1_2_4_en,
    output[1:0] io_VwirePorts_1_2_4_out,
    input [1:0] io_VwirePorts_1_2_3_in,
    input  io_VwirePorts_1_2_3_en,
    output[1:0] io_VwirePorts_1_2_3_out,
    input [1:0] io_VwirePorts_1_2_2_in,
    input  io_VwirePorts_1_2_2_en,
    output[1:0] io_VwirePorts_1_2_2_out,
    input [1:0] io_VwirePorts_1_2_1_in,
    input  io_VwirePorts_1_2_1_en,
    output[1:0] io_VwirePorts_1_2_1_out,
    input [1:0] io_VwirePorts_1_2_0_in,
    input  io_VwirePorts_1_2_0_en,
    output[1:0] io_VwirePorts_1_2_0_out,
    input [1:0] io_VwirePorts_1_1_15_in,
    input  io_VwirePorts_1_1_15_en,
    output[1:0] io_VwirePorts_1_1_15_out,
    input [1:0] io_VwirePorts_1_1_14_in,
    input  io_VwirePorts_1_1_14_en,
    output[1:0] io_VwirePorts_1_1_14_out,
    input [1:0] io_VwirePorts_1_1_13_in,
    input  io_VwirePorts_1_1_13_en,
    output[1:0] io_VwirePorts_1_1_13_out,
    input [1:0] io_VwirePorts_1_1_12_in,
    input  io_VwirePorts_1_1_12_en,
    output[1:0] io_VwirePorts_1_1_12_out,
    input [1:0] io_VwirePorts_1_1_11_in,
    input  io_VwirePorts_1_1_11_en,
    output[1:0] io_VwirePorts_1_1_11_out,
    input [1:0] io_VwirePorts_1_1_10_in,
    input  io_VwirePorts_1_1_10_en,
    output[1:0] io_VwirePorts_1_1_10_out,
    input [1:0] io_VwirePorts_1_1_9_in,
    input  io_VwirePorts_1_1_9_en,
    output[1:0] io_VwirePorts_1_1_9_out,
    input [1:0] io_VwirePorts_1_1_8_in,
    input  io_VwirePorts_1_1_8_en,
    output[1:0] io_VwirePorts_1_1_8_out,
    input [1:0] io_VwirePorts_1_1_7_in,
    input  io_VwirePorts_1_1_7_en,
    output[1:0] io_VwirePorts_1_1_7_out,
    input [1:0] io_VwirePorts_1_1_6_in,
    input  io_VwirePorts_1_1_6_en,
    output[1:0] io_VwirePorts_1_1_6_out,
    input [1:0] io_VwirePorts_1_1_5_in,
    input  io_VwirePorts_1_1_5_en,
    output[1:0] io_VwirePorts_1_1_5_out,
    input [1:0] io_VwirePorts_1_1_4_in,
    input  io_VwirePorts_1_1_4_en,
    output[1:0] io_VwirePorts_1_1_4_out,
    input [1:0] io_VwirePorts_1_1_3_in,
    input  io_VwirePorts_1_1_3_en,
    output[1:0] io_VwirePorts_1_1_3_out,
    input [1:0] io_VwirePorts_1_1_2_in,
    input  io_VwirePorts_1_1_2_en,
    output[1:0] io_VwirePorts_1_1_2_out,
    input [1:0] io_VwirePorts_1_1_1_in,
    input  io_VwirePorts_1_1_1_en,
    output[1:0] io_VwirePorts_1_1_1_out,
    input [1:0] io_VwirePorts_1_1_0_in,
    input  io_VwirePorts_1_1_0_en,
    output[1:0] io_VwirePorts_1_1_0_out,
    input [1:0] io_VwirePorts_1_0_15_in,
    input  io_VwirePorts_1_0_15_en,
    output[1:0] io_VwirePorts_1_0_15_out,
    input [1:0] io_VwirePorts_1_0_14_in,
    input  io_VwirePorts_1_0_14_en,
    output[1:0] io_VwirePorts_1_0_14_out,
    input [1:0] io_VwirePorts_1_0_13_in,
    input  io_VwirePorts_1_0_13_en,
    output[1:0] io_VwirePorts_1_0_13_out,
    input [1:0] io_VwirePorts_1_0_12_in,
    input  io_VwirePorts_1_0_12_en,
    output[1:0] io_VwirePorts_1_0_12_out,
    input [1:0] io_VwirePorts_1_0_11_in,
    input  io_VwirePorts_1_0_11_en,
    output[1:0] io_VwirePorts_1_0_11_out,
    input [1:0] io_VwirePorts_1_0_10_in,
    input  io_VwirePorts_1_0_10_en,
    output[1:0] io_VwirePorts_1_0_10_out,
    input [1:0] io_VwirePorts_1_0_9_in,
    input  io_VwirePorts_1_0_9_en,
    output[1:0] io_VwirePorts_1_0_9_out,
    input [1:0] io_VwirePorts_1_0_8_in,
    input  io_VwirePorts_1_0_8_en,
    output[1:0] io_VwirePorts_1_0_8_out,
    input [1:0] io_VwirePorts_1_0_7_in,
    input  io_VwirePorts_1_0_7_en,
    output[1:0] io_VwirePorts_1_0_7_out,
    input [1:0] io_VwirePorts_1_0_6_in,
    input  io_VwirePorts_1_0_6_en,
    output[1:0] io_VwirePorts_1_0_6_out,
    input [1:0] io_VwirePorts_1_0_5_in,
    input  io_VwirePorts_1_0_5_en,
    output[1:0] io_VwirePorts_1_0_5_out,
    input [1:0] io_VwirePorts_1_0_4_in,
    input  io_VwirePorts_1_0_4_en,
    output[1:0] io_VwirePorts_1_0_4_out,
    input [1:0] io_VwirePorts_1_0_3_in,
    input  io_VwirePorts_1_0_3_en,
    output[1:0] io_VwirePorts_1_0_3_out,
    input [1:0] io_VwirePorts_1_0_2_in,
    input  io_VwirePorts_1_0_2_en,
    output[1:0] io_VwirePorts_1_0_2_out,
    input [1:0] io_VwirePorts_1_0_1_in,
    input  io_VwirePorts_1_0_1_en,
    output[1:0] io_VwirePorts_1_0_1_out,
    input [1:0] io_VwirePorts_1_0_0_in,
    input  io_VwirePorts_1_0_0_en,
    output[1:0] io_VwirePorts_1_0_0_out,
    input [1:0] io_VwirePorts_0_22_15_in,
    input  io_VwirePorts_0_22_15_en,
    output[1:0] io_VwirePorts_0_22_15_out,
    input [1:0] io_VwirePorts_0_22_14_in,
    input  io_VwirePorts_0_22_14_en,
    output[1:0] io_VwirePorts_0_22_14_out,
    input [1:0] io_VwirePorts_0_22_13_in,
    input  io_VwirePorts_0_22_13_en,
    output[1:0] io_VwirePorts_0_22_13_out,
    input [1:0] io_VwirePorts_0_22_12_in,
    input  io_VwirePorts_0_22_12_en,
    output[1:0] io_VwirePorts_0_22_12_out,
    input [1:0] io_VwirePorts_0_22_11_in,
    input  io_VwirePorts_0_22_11_en,
    output[1:0] io_VwirePorts_0_22_11_out,
    input [1:0] io_VwirePorts_0_22_10_in,
    input  io_VwirePorts_0_22_10_en,
    output[1:0] io_VwirePorts_0_22_10_out,
    input [1:0] io_VwirePorts_0_22_9_in,
    input  io_VwirePorts_0_22_9_en,
    output[1:0] io_VwirePorts_0_22_9_out,
    input [1:0] io_VwirePorts_0_22_8_in,
    input  io_VwirePorts_0_22_8_en,
    output[1:0] io_VwirePorts_0_22_8_out,
    input [1:0] io_VwirePorts_0_22_7_in,
    input  io_VwirePorts_0_22_7_en,
    output[1:0] io_VwirePorts_0_22_7_out,
    input [1:0] io_VwirePorts_0_22_6_in,
    input  io_VwirePorts_0_22_6_en,
    output[1:0] io_VwirePorts_0_22_6_out,
    input [1:0] io_VwirePorts_0_22_5_in,
    input  io_VwirePorts_0_22_5_en,
    output[1:0] io_VwirePorts_0_22_5_out,
    input [1:0] io_VwirePorts_0_22_4_in,
    input  io_VwirePorts_0_22_4_en,
    output[1:0] io_VwirePorts_0_22_4_out,
    input [1:0] io_VwirePorts_0_22_3_in,
    input  io_VwirePorts_0_22_3_en,
    output[1:0] io_VwirePorts_0_22_3_out,
    input [1:0] io_VwirePorts_0_22_2_in,
    input  io_VwirePorts_0_22_2_en,
    output[1:0] io_VwirePorts_0_22_2_out,
    input [1:0] io_VwirePorts_0_22_1_in,
    input  io_VwirePorts_0_22_1_en,
    output[1:0] io_VwirePorts_0_22_1_out,
    input [1:0] io_VwirePorts_0_22_0_in,
    input  io_VwirePorts_0_22_0_en,
    output[1:0] io_VwirePorts_0_22_0_out,
    input [1:0] io_VwirePorts_0_21_15_in,
    input  io_VwirePorts_0_21_15_en,
    output[1:0] io_VwirePorts_0_21_15_out,
    input [1:0] io_VwirePorts_0_21_14_in,
    input  io_VwirePorts_0_21_14_en,
    output[1:0] io_VwirePorts_0_21_14_out,
    input [1:0] io_VwirePorts_0_21_13_in,
    input  io_VwirePorts_0_21_13_en,
    output[1:0] io_VwirePorts_0_21_13_out,
    input [1:0] io_VwirePorts_0_21_12_in,
    input  io_VwirePorts_0_21_12_en,
    output[1:0] io_VwirePorts_0_21_12_out,
    input [1:0] io_VwirePorts_0_21_11_in,
    input  io_VwirePorts_0_21_11_en,
    output[1:0] io_VwirePorts_0_21_11_out,
    input [1:0] io_VwirePorts_0_21_10_in,
    input  io_VwirePorts_0_21_10_en,
    output[1:0] io_VwirePorts_0_21_10_out,
    input [1:0] io_VwirePorts_0_21_9_in,
    input  io_VwirePorts_0_21_9_en,
    output[1:0] io_VwirePorts_0_21_9_out,
    input [1:0] io_VwirePorts_0_21_8_in,
    input  io_VwirePorts_0_21_8_en,
    output[1:0] io_VwirePorts_0_21_8_out,
    input [1:0] io_VwirePorts_0_21_7_in,
    input  io_VwirePorts_0_21_7_en,
    output[1:0] io_VwirePorts_0_21_7_out,
    input [1:0] io_VwirePorts_0_21_6_in,
    input  io_VwirePorts_0_21_6_en,
    output[1:0] io_VwirePorts_0_21_6_out,
    input [1:0] io_VwirePorts_0_21_5_in,
    input  io_VwirePorts_0_21_5_en,
    output[1:0] io_VwirePorts_0_21_5_out,
    input [1:0] io_VwirePorts_0_21_4_in,
    input  io_VwirePorts_0_21_4_en,
    output[1:0] io_VwirePorts_0_21_4_out,
    input [1:0] io_VwirePorts_0_21_3_in,
    input  io_VwirePorts_0_21_3_en,
    output[1:0] io_VwirePorts_0_21_3_out,
    input [1:0] io_VwirePorts_0_21_2_in,
    input  io_VwirePorts_0_21_2_en,
    output[1:0] io_VwirePorts_0_21_2_out,
    input [1:0] io_VwirePorts_0_21_1_in,
    input  io_VwirePorts_0_21_1_en,
    output[1:0] io_VwirePorts_0_21_1_out,
    input [1:0] io_VwirePorts_0_21_0_in,
    input  io_VwirePorts_0_21_0_en,
    output[1:0] io_VwirePorts_0_21_0_out,
    input [1:0] io_VwirePorts_0_20_15_in,
    input  io_VwirePorts_0_20_15_en,
    output[1:0] io_VwirePorts_0_20_15_out,
    input [1:0] io_VwirePorts_0_20_14_in,
    input  io_VwirePorts_0_20_14_en,
    output[1:0] io_VwirePorts_0_20_14_out,
    input [1:0] io_VwirePorts_0_20_13_in,
    input  io_VwirePorts_0_20_13_en,
    output[1:0] io_VwirePorts_0_20_13_out,
    input [1:0] io_VwirePorts_0_20_12_in,
    input  io_VwirePorts_0_20_12_en,
    output[1:0] io_VwirePorts_0_20_12_out,
    input [1:0] io_VwirePorts_0_20_11_in,
    input  io_VwirePorts_0_20_11_en,
    output[1:0] io_VwirePorts_0_20_11_out,
    input [1:0] io_VwirePorts_0_20_10_in,
    input  io_VwirePorts_0_20_10_en,
    output[1:0] io_VwirePorts_0_20_10_out,
    input [1:0] io_VwirePorts_0_20_9_in,
    input  io_VwirePorts_0_20_9_en,
    output[1:0] io_VwirePorts_0_20_9_out,
    input [1:0] io_VwirePorts_0_20_8_in,
    input  io_VwirePorts_0_20_8_en,
    output[1:0] io_VwirePorts_0_20_8_out,
    input [1:0] io_VwirePorts_0_20_7_in,
    input  io_VwirePorts_0_20_7_en,
    output[1:0] io_VwirePorts_0_20_7_out,
    input [1:0] io_VwirePorts_0_20_6_in,
    input  io_VwirePorts_0_20_6_en,
    output[1:0] io_VwirePorts_0_20_6_out,
    input [1:0] io_VwirePorts_0_20_5_in,
    input  io_VwirePorts_0_20_5_en,
    output[1:0] io_VwirePorts_0_20_5_out,
    input [1:0] io_VwirePorts_0_20_4_in,
    input  io_VwirePorts_0_20_4_en,
    output[1:0] io_VwirePorts_0_20_4_out,
    input [1:0] io_VwirePorts_0_20_3_in,
    input  io_VwirePorts_0_20_3_en,
    output[1:0] io_VwirePorts_0_20_3_out,
    input [1:0] io_VwirePorts_0_20_2_in,
    input  io_VwirePorts_0_20_2_en,
    output[1:0] io_VwirePorts_0_20_2_out,
    input [1:0] io_VwirePorts_0_20_1_in,
    input  io_VwirePorts_0_20_1_en,
    output[1:0] io_VwirePorts_0_20_1_out,
    input [1:0] io_VwirePorts_0_20_0_in,
    input  io_VwirePorts_0_20_0_en,
    output[1:0] io_VwirePorts_0_20_0_out,
    input [1:0] io_VwirePorts_0_19_15_in,
    input  io_VwirePorts_0_19_15_en,
    output[1:0] io_VwirePorts_0_19_15_out,
    input [1:0] io_VwirePorts_0_19_14_in,
    input  io_VwirePorts_0_19_14_en,
    output[1:0] io_VwirePorts_0_19_14_out,
    input [1:0] io_VwirePorts_0_19_13_in,
    input  io_VwirePorts_0_19_13_en,
    output[1:0] io_VwirePorts_0_19_13_out,
    input [1:0] io_VwirePorts_0_19_12_in,
    input  io_VwirePorts_0_19_12_en,
    output[1:0] io_VwirePorts_0_19_12_out,
    input [1:0] io_VwirePorts_0_19_11_in,
    input  io_VwirePorts_0_19_11_en,
    output[1:0] io_VwirePorts_0_19_11_out,
    input [1:0] io_VwirePorts_0_19_10_in,
    input  io_VwirePorts_0_19_10_en,
    output[1:0] io_VwirePorts_0_19_10_out,
    input [1:0] io_VwirePorts_0_19_9_in,
    input  io_VwirePorts_0_19_9_en,
    output[1:0] io_VwirePorts_0_19_9_out,
    input [1:0] io_VwirePorts_0_19_8_in,
    input  io_VwirePorts_0_19_8_en,
    output[1:0] io_VwirePorts_0_19_8_out,
    input [1:0] io_VwirePorts_0_19_7_in,
    input  io_VwirePorts_0_19_7_en,
    output[1:0] io_VwirePorts_0_19_7_out,
    input [1:0] io_VwirePorts_0_19_6_in,
    input  io_VwirePorts_0_19_6_en,
    output[1:0] io_VwirePorts_0_19_6_out,
    input [1:0] io_VwirePorts_0_19_5_in,
    input  io_VwirePorts_0_19_5_en,
    output[1:0] io_VwirePorts_0_19_5_out,
    input [1:0] io_VwirePorts_0_19_4_in,
    input  io_VwirePorts_0_19_4_en,
    output[1:0] io_VwirePorts_0_19_4_out,
    input [1:0] io_VwirePorts_0_19_3_in,
    input  io_VwirePorts_0_19_3_en,
    output[1:0] io_VwirePorts_0_19_3_out,
    input [1:0] io_VwirePorts_0_19_2_in,
    input  io_VwirePorts_0_19_2_en,
    output[1:0] io_VwirePorts_0_19_2_out,
    input [1:0] io_VwirePorts_0_19_1_in,
    input  io_VwirePorts_0_19_1_en,
    output[1:0] io_VwirePorts_0_19_1_out,
    input [1:0] io_VwirePorts_0_19_0_in,
    input  io_VwirePorts_0_19_0_en,
    output[1:0] io_VwirePorts_0_19_0_out,
    input [1:0] io_VwirePorts_0_18_15_in,
    input  io_VwirePorts_0_18_15_en,
    output[1:0] io_VwirePorts_0_18_15_out,
    input [1:0] io_VwirePorts_0_18_14_in,
    input  io_VwirePorts_0_18_14_en,
    output[1:0] io_VwirePorts_0_18_14_out,
    input [1:0] io_VwirePorts_0_18_13_in,
    input  io_VwirePorts_0_18_13_en,
    output[1:0] io_VwirePorts_0_18_13_out,
    input [1:0] io_VwirePorts_0_18_12_in,
    input  io_VwirePorts_0_18_12_en,
    output[1:0] io_VwirePorts_0_18_12_out,
    input [1:0] io_VwirePorts_0_18_11_in,
    input  io_VwirePorts_0_18_11_en,
    output[1:0] io_VwirePorts_0_18_11_out,
    input [1:0] io_VwirePorts_0_18_10_in,
    input  io_VwirePorts_0_18_10_en,
    output[1:0] io_VwirePorts_0_18_10_out,
    input [1:0] io_VwirePorts_0_18_9_in,
    input  io_VwirePorts_0_18_9_en,
    output[1:0] io_VwirePorts_0_18_9_out,
    input [1:0] io_VwirePorts_0_18_8_in,
    input  io_VwirePorts_0_18_8_en,
    output[1:0] io_VwirePorts_0_18_8_out,
    input [1:0] io_VwirePorts_0_18_7_in,
    input  io_VwirePorts_0_18_7_en,
    output[1:0] io_VwirePorts_0_18_7_out,
    input [1:0] io_VwirePorts_0_18_6_in,
    input  io_VwirePorts_0_18_6_en,
    output[1:0] io_VwirePorts_0_18_6_out,
    input [1:0] io_VwirePorts_0_18_5_in,
    input  io_VwirePorts_0_18_5_en,
    output[1:0] io_VwirePorts_0_18_5_out,
    input [1:0] io_VwirePorts_0_18_4_in,
    input  io_VwirePorts_0_18_4_en,
    output[1:0] io_VwirePorts_0_18_4_out,
    input [1:0] io_VwirePorts_0_18_3_in,
    input  io_VwirePorts_0_18_3_en,
    output[1:0] io_VwirePorts_0_18_3_out,
    input [1:0] io_VwirePorts_0_18_2_in,
    input  io_VwirePorts_0_18_2_en,
    output[1:0] io_VwirePorts_0_18_2_out,
    input [1:0] io_VwirePorts_0_18_1_in,
    input  io_VwirePorts_0_18_1_en,
    output[1:0] io_VwirePorts_0_18_1_out,
    input [1:0] io_VwirePorts_0_18_0_in,
    input  io_VwirePorts_0_18_0_en,
    output[1:0] io_VwirePorts_0_18_0_out,
    input [1:0] io_VwirePorts_0_17_15_in,
    input  io_VwirePorts_0_17_15_en,
    output[1:0] io_VwirePorts_0_17_15_out,
    input [1:0] io_VwirePorts_0_17_14_in,
    input  io_VwirePorts_0_17_14_en,
    output[1:0] io_VwirePorts_0_17_14_out,
    input [1:0] io_VwirePorts_0_17_13_in,
    input  io_VwirePorts_0_17_13_en,
    output[1:0] io_VwirePorts_0_17_13_out,
    input [1:0] io_VwirePorts_0_17_12_in,
    input  io_VwirePorts_0_17_12_en,
    output[1:0] io_VwirePorts_0_17_12_out,
    input [1:0] io_VwirePorts_0_17_11_in,
    input  io_VwirePorts_0_17_11_en,
    output[1:0] io_VwirePorts_0_17_11_out,
    input [1:0] io_VwirePorts_0_17_10_in,
    input  io_VwirePorts_0_17_10_en,
    output[1:0] io_VwirePorts_0_17_10_out,
    input [1:0] io_VwirePorts_0_17_9_in,
    input  io_VwirePorts_0_17_9_en,
    output[1:0] io_VwirePorts_0_17_9_out,
    input [1:0] io_VwirePorts_0_17_8_in,
    input  io_VwirePorts_0_17_8_en,
    output[1:0] io_VwirePorts_0_17_8_out,
    input [1:0] io_VwirePorts_0_17_7_in,
    input  io_VwirePorts_0_17_7_en,
    output[1:0] io_VwirePorts_0_17_7_out,
    input [1:0] io_VwirePorts_0_17_6_in,
    input  io_VwirePorts_0_17_6_en,
    output[1:0] io_VwirePorts_0_17_6_out,
    input [1:0] io_VwirePorts_0_17_5_in,
    input  io_VwirePorts_0_17_5_en,
    output[1:0] io_VwirePorts_0_17_5_out,
    input [1:0] io_VwirePorts_0_17_4_in,
    input  io_VwirePorts_0_17_4_en,
    output[1:0] io_VwirePorts_0_17_4_out,
    input [1:0] io_VwirePorts_0_17_3_in,
    input  io_VwirePorts_0_17_3_en,
    output[1:0] io_VwirePorts_0_17_3_out,
    input [1:0] io_VwirePorts_0_17_2_in,
    input  io_VwirePorts_0_17_2_en,
    output[1:0] io_VwirePorts_0_17_2_out,
    input [1:0] io_VwirePorts_0_17_1_in,
    input  io_VwirePorts_0_17_1_en,
    output[1:0] io_VwirePorts_0_17_1_out,
    input [1:0] io_VwirePorts_0_17_0_in,
    input  io_VwirePorts_0_17_0_en,
    output[1:0] io_VwirePorts_0_17_0_out,
    input [1:0] io_VwirePorts_0_16_15_in,
    input  io_VwirePorts_0_16_15_en,
    output[1:0] io_VwirePorts_0_16_15_out,
    input [1:0] io_VwirePorts_0_16_14_in,
    input  io_VwirePorts_0_16_14_en,
    output[1:0] io_VwirePorts_0_16_14_out,
    input [1:0] io_VwirePorts_0_16_13_in,
    input  io_VwirePorts_0_16_13_en,
    output[1:0] io_VwirePorts_0_16_13_out,
    input [1:0] io_VwirePorts_0_16_12_in,
    input  io_VwirePorts_0_16_12_en,
    output[1:0] io_VwirePorts_0_16_12_out,
    input [1:0] io_VwirePorts_0_16_11_in,
    input  io_VwirePorts_0_16_11_en,
    output[1:0] io_VwirePorts_0_16_11_out,
    input [1:0] io_VwirePorts_0_16_10_in,
    input  io_VwirePorts_0_16_10_en,
    output[1:0] io_VwirePorts_0_16_10_out,
    input [1:0] io_VwirePorts_0_16_9_in,
    input  io_VwirePorts_0_16_9_en,
    output[1:0] io_VwirePorts_0_16_9_out,
    input [1:0] io_VwirePorts_0_16_8_in,
    input  io_VwirePorts_0_16_8_en,
    output[1:0] io_VwirePorts_0_16_8_out,
    input [1:0] io_VwirePorts_0_16_7_in,
    input  io_VwirePorts_0_16_7_en,
    output[1:0] io_VwirePorts_0_16_7_out,
    input [1:0] io_VwirePorts_0_16_6_in,
    input  io_VwirePorts_0_16_6_en,
    output[1:0] io_VwirePorts_0_16_6_out,
    input [1:0] io_VwirePorts_0_16_5_in,
    input  io_VwirePorts_0_16_5_en,
    output[1:0] io_VwirePorts_0_16_5_out,
    input [1:0] io_VwirePorts_0_16_4_in,
    input  io_VwirePorts_0_16_4_en,
    output[1:0] io_VwirePorts_0_16_4_out,
    input [1:0] io_VwirePorts_0_16_3_in,
    input  io_VwirePorts_0_16_3_en,
    output[1:0] io_VwirePorts_0_16_3_out,
    input [1:0] io_VwirePorts_0_16_2_in,
    input  io_VwirePorts_0_16_2_en,
    output[1:0] io_VwirePorts_0_16_2_out,
    input [1:0] io_VwirePorts_0_16_1_in,
    input  io_VwirePorts_0_16_1_en,
    output[1:0] io_VwirePorts_0_16_1_out,
    input [1:0] io_VwirePorts_0_16_0_in,
    input  io_VwirePorts_0_16_0_en,
    output[1:0] io_VwirePorts_0_16_0_out,
    input [1:0] io_VwirePorts_0_15_15_in,
    input  io_VwirePorts_0_15_15_en,
    output[1:0] io_VwirePorts_0_15_15_out,
    input [1:0] io_VwirePorts_0_15_14_in,
    input  io_VwirePorts_0_15_14_en,
    output[1:0] io_VwirePorts_0_15_14_out,
    input [1:0] io_VwirePorts_0_15_13_in,
    input  io_VwirePorts_0_15_13_en,
    output[1:0] io_VwirePorts_0_15_13_out,
    input [1:0] io_VwirePorts_0_15_12_in,
    input  io_VwirePorts_0_15_12_en,
    output[1:0] io_VwirePorts_0_15_12_out,
    input [1:0] io_VwirePorts_0_15_11_in,
    input  io_VwirePorts_0_15_11_en,
    output[1:0] io_VwirePorts_0_15_11_out,
    input [1:0] io_VwirePorts_0_15_10_in,
    input  io_VwirePorts_0_15_10_en,
    output[1:0] io_VwirePorts_0_15_10_out,
    input [1:0] io_VwirePorts_0_15_9_in,
    input  io_VwirePorts_0_15_9_en,
    output[1:0] io_VwirePorts_0_15_9_out,
    input [1:0] io_VwirePorts_0_15_8_in,
    input  io_VwirePorts_0_15_8_en,
    output[1:0] io_VwirePorts_0_15_8_out,
    input [1:0] io_VwirePorts_0_15_7_in,
    input  io_VwirePorts_0_15_7_en,
    output[1:0] io_VwirePorts_0_15_7_out,
    input [1:0] io_VwirePorts_0_15_6_in,
    input  io_VwirePorts_0_15_6_en,
    output[1:0] io_VwirePorts_0_15_6_out,
    input [1:0] io_VwirePorts_0_15_5_in,
    input  io_VwirePorts_0_15_5_en,
    output[1:0] io_VwirePorts_0_15_5_out,
    input [1:0] io_VwirePorts_0_15_4_in,
    input  io_VwirePorts_0_15_4_en,
    output[1:0] io_VwirePorts_0_15_4_out,
    input [1:0] io_VwirePorts_0_15_3_in,
    input  io_VwirePorts_0_15_3_en,
    output[1:0] io_VwirePorts_0_15_3_out,
    input [1:0] io_VwirePorts_0_15_2_in,
    input  io_VwirePorts_0_15_2_en,
    output[1:0] io_VwirePorts_0_15_2_out,
    input [1:0] io_VwirePorts_0_15_1_in,
    input  io_VwirePorts_0_15_1_en,
    output[1:0] io_VwirePorts_0_15_1_out,
    input [1:0] io_VwirePorts_0_15_0_in,
    input  io_VwirePorts_0_15_0_en,
    output[1:0] io_VwirePorts_0_15_0_out,
    input [1:0] io_VwirePorts_0_14_15_in,
    input  io_VwirePorts_0_14_15_en,
    output[1:0] io_VwirePorts_0_14_15_out,
    input [1:0] io_VwirePorts_0_14_14_in,
    input  io_VwirePorts_0_14_14_en,
    output[1:0] io_VwirePorts_0_14_14_out,
    input [1:0] io_VwirePorts_0_14_13_in,
    input  io_VwirePorts_0_14_13_en,
    output[1:0] io_VwirePorts_0_14_13_out,
    input [1:0] io_VwirePorts_0_14_12_in,
    input  io_VwirePorts_0_14_12_en,
    output[1:0] io_VwirePorts_0_14_12_out,
    input [1:0] io_VwirePorts_0_14_11_in,
    input  io_VwirePorts_0_14_11_en,
    output[1:0] io_VwirePorts_0_14_11_out,
    input [1:0] io_VwirePorts_0_14_10_in,
    input  io_VwirePorts_0_14_10_en,
    output[1:0] io_VwirePorts_0_14_10_out,
    input [1:0] io_VwirePorts_0_14_9_in,
    input  io_VwirePorts_0_14_9_en,
    output[1:0] io_VwirePorts_0_14_9_out,
    input [1:0] io_VwirePorts_0_14_8_in,
    input  io_VwirePorts_0_14_8_en,
    output[1:0] io_VwirePorts_0_14_8_out,
    input [1:0] io_VwirePorts_0_14_7_in,
    input  io_VwirePorts_0_14_7_en,
    output[1:0] io_VwirePorts_0_14_7_out,
    input [1:0] io_VwirePorts_0_14_6_in,
    input  io_VwirePorts_0_14_6_en,
    output[1:0] io_VwirePorts_0_14_6_out,
    input [1:0] io_VwirePorts_0_14_5_in,
    input  io_VwirePorts_0_14_5_en,
    output[1:0] io_VwirePorts_0_14_5_out,
    input [1:0] io_VwirePorts_0_14_4_in,
    input  io_VwirePorts_0_14_4_en,
    output[1:0] io_VwirePorts_0_14_4_out,
    input [1:0] io_VwirePorts_0_14_3_in,
    input  io_VwirePorts_0_14_3_en,
    output[1:0] io_VwirePorts_0_14_3_out,
    input [1:0] io_VwirePorts_0_14_2_in,
    input  io_VwirePorts_0_14_2_en,
    output[1:0] io_VwirePorts_0_14_2_out,
    input [1:0] io_VwirePorts_0_14_1_in,
    input  io_VwirePorts_0_14_1_en,
    output[1:0] io_VwirePorts_0_14_1_out,
    input [1:0] io_VwirePorts_0_14_0_in,
    input  io_VwirePorts_0_14_0_en,
    output[1:0] io_VwirePorts_0_14_0_out,
    input [1:0] io_VwirePorts_0_13_15_in,
    input  io_VwirePorts_0_13_15_en,
    output[1:0] io_VwirePorts_0_13_15_out,
    input [1:0] io_VwirePorts_0_13_14_in,
    input  io_VwirePorts_0_13_14_en,
    output[1:0] io_VwirePorts_0_13_14_out,
    input [1:0] io_VwirePorts_0_13_13_in,
    input  io_VwirePorts_0_13_13_en,
    output[1:0] io_VwirePorts_0_13_13_out,
    input [1:0] io_VwirePorts_0_13_12_in,
    input  io_VwirePorts_0_13_12_en,
    output[1:0] io_VwirePorts_0_13_12_out,
    input [1:0] io_VwirePorts_0_13_11_in,
    input  io_VwirePorts_0_13_11_en,
    output[1:0] io_VwirePorts_0_13_11_out,
    input [1:0] io_VwirePorts_0_13_10_in,
    input  io_VwirePorts_0_13_10_en,
    output[1:0] io_VwirePorts_0_13_10_out,
    input [1:0] io_VwirePorts_0_13_9_in,
    input  io_VwirePorts_0_13_9_en,
    output[1:0] io_VwirePorts_0_13_9_out,
    input [1:0] io_VwirePorts_0_13_8_in,
    input  io_VwirePorts_0_13_8_en,
    output[1:0] io_VwirePorts_0_13_8_out,
    input [1:0] io_VwirePorts_0_13_7_in,
    input  io_VwirePorts_0_13_7_en,
    output[1:0] io_VwirePorts_0_13_7_out,
    input [1:0] io_VwirePorts_0_13_6_in,
    input  io_VwirePorts_0_13_6_en,
    output[1:0] io_VwirePorts_0_13_6_out,
    input [1:0] io_VwirePorts_0_13_5_in,
    input  io_VwirePorts_0_13_5_en,
    output[1:0] io_VwirePorts_0_13_5_out,
    input [1:0] io_VwirePorts_0_13_4_in,
    input  io_VwirePorts_0_13_4_en,
    output[1:0] io_VwirePorts_0_13_4_out,
    input [1:0] io_VwirePorts_0_13_3_in,
    input  io_VwirePorts_0_13_3_en,
    output[1:0] io_VwirePorts_0_13_3_out,
    input [1:0] io_VwirePorts_0_13_2_in,
    input  io_VwirePorts_0_13_2_en,
    output[1:0] io_VwirePorts_0_13_2_out,
    input [1:0] io_VwirePorts_0_13_1_in,
    input  io_VwirePorts_0_13_1_en,
    output[1:0] io_VwirePorts_0_13_1_out,
    input [1:0] io_VwirePorts_0_13_0_in,
    input  io_VwirePorts_0_13_0_en,
    output[1:0] io_VwirePorts_0_13_0_out,
    input [1:0] io_VwirePorts_0_12_15_in,
    input  io_VwirePorts_0_12_15_en,
    output[1:0] io_VwirePorts_0_12_15_out,
    input [1:0] io_VwirePorts_0_12_14_in,
    input  io_VwirePorts_0_12_14_en,
    output[1:0] io_VwirePorts_0_12_14_out,
    input [1:0] io_VwirePorts_0_12_13_in,
    input  io_VwirePorts_0_12_13_en,
    output[1:0] io_VwirePorts_0_12_13_out,
    input [1:0] io_VwirePorts_0_12_12_in,
    input  io_VwirePorts_0_12_12_en,
    output[1:0] io_VwirePorts_0_12_12_out,
    input [1:0] io_VwirePorts_0_12_11_in,
    input  io_VwirePorts_0_12_11_en,
    output[1:0] io_VwirePorts_0_12_11_out,
    input [1:0] io_VwirePorts_0_12_10_in,
    input  io_VwirePorts_0_12_10_en,
    output[1:0] io_VwirePorts_0_12_10_out,
    input [1:0] io_VwirePorts_0_12_9_in,
    input  io_VwirePorts_0_12_9_en,
    output[1:0] io_VwirePorts_0_12_9_out,
    input [1:0] io_VwirePorts_0_12_8_in,
    input  io_VwirePorts_0_12_8_en,
    output[1:0] io_VwirePorts_0_12_8_out,
    input [1:0] io_VwirePorts_0_12_7_in,
    input  io_VwirePorts_0_12_7_en,
    output[1:0] io_VwirePorts_0_12_7_out,
    input [1:0] io_VwirePorts_0_12_6_in,
    input  io_VwirePorts_0_12_6_en,
    output[1:0] io_VwirePorts_0_12_6_out,
    input [1:0] io_VwirePorts_0_12_5_in,
    input  io_VwirePorts_0_12_5_en,
    output[1:0] io_VwirePorts_0_12_5_out,
    input [1:0] io_VwirePorts_0_12_4_in,
    input  io_VwirePorts_0_12_4_en,
    output[1:0] io_VwirePorts_0_12_4_out,
    input [1:0] io_VwirePorts_0_12_3_in,
    input  io_VwirePorts_0_12_3_en,
    output[1:0] io_VwirePorts_0_12_3_out,
    input [1:0] io_VwirePorts_0_12_2_in,
    input  io_VwirePorts_0_12_2_en,
    output[1:0] io_VwirePorts_0_12_2_out,
    input [1:0] io_VwirePorts_0_12_1_in,
    input  io_VwirePorts_0_12_1_en,
    output[1:0] io_VwirePorts_0_12_1_out,
    input [1:0] io_VwirePorts_0_12_0_in,
    input  io_VwirePorts_0_12_0_en,
    output[1:0] io_VwirePorts_0_12_0_out,
    input [1:0] io_VwirePorts_0_11_15_in,
    input  io_VwirePorts_0_11_15_en,
    output[1:0] io_VwirePorts_0_11_15_out,
    input [1:0] io_VwirePorts_0_11_14_in,
    input  io_VwirePorts_0_11_14_en,
    output[1:0] io_VwirePorts_0_11_14_out,
    input [1:0] io_VwirePorts_0_11_13_in,
    input  io_VwirePorts_0_11_13_en,
    output[1:0] io_VwirePorts_0_11_13_out,
    input [1:0] io_VwirePorts_0_11_12_in,
    input  io_VwirePorts_0_11_12_en,
    output[1:0] io_VwirePorts_0_11_12_out,
    input [1:0] io_VwirePorts_0_11_11_in,
    input  io_VwirePorts_0_11_11_en,
    output[1:0] io_VwirePorts_0_11_11_out,
    input [1:0] io_VwirePorts_0_11_10_in,
    input  io_VwirePorts_0_11_10_en,
    output[1:0] io_VwirePorts_0_11_10_out,
    input [1:0] io_VwirePorts_0_11_9_in,
    input  io_VwirePorts_0_11_9_en,
    output[1:0] io_VwirePorts_0_11_9_out,
    input [1:0] io_VwirePorts_0_11_8_in,
    input  io_VwirePorts_0_11_8_en,
    output[1:0] io_VwirePorts_0_11_8_out,
    input [1:0] io_VwirePorts_0_11_7_in,
    input  io_VwirePorts_0_11_7_en,
    output[1:0] io_VwirePorts_0_11_7_out,
    input [1:0] io_VwirePorts_0_11_6_in,
    input  io_VwirePorts_0_11_6_en,
    output[1:0] io_VwirePorts_0_11_6_out,
    input [1:0] io_VwirePorts_0_11_5_in,
    input  io_VwirePorts_0_11_5_en,
    output[1:0] io_VwirePorts_0_11_5_out,
    input [1:0] io_VwirePorts_0_11_4_in,
    input  io_VwirePorts_0_11_4_en,
    output[1:0] io_VwirePorts_0_11_4_out,
    input [1:0] io_VwirePorts_0_11_3_in,
    input  io_VwirePorts_0_11_3_en,
    output[1:0] io_VwirePorts_0_11_3_out,
    input [1:0] io_VwirePorts_0_11_2_in,
    input  io_VwirePorts_0_11_2_en,
    output[1:0] io_VwirePorts_0_11_2_out,
    input [1:0] io_VwirePorts_0_11_1_in,
    input  io_VwirePorts_0_11_1_en,
    output[1:0] io_VwirePorts_0_11_1_out,
    input [1:0] io_VwirePorts_0_11_0_in,
    input  io_VwirePorts_0_11_0_en,
    output[1:0] io_VwirePorts_0_11_0_out,
    input [1:0] io_VwirePorts_0_10_15_in,
    input  io_VwirePorts_0_10_15_en,
    output[1:0] io_VwirePorts_0_10_15_out,
    input [1:0] io_VwirePorts_0_10_14_in,
    input  io_VwirePorts_0_10_14_en,
    output[1:0] io_VwirePorts_0_10_14_out,
    input [1:0] io_VwirePorts_0_10_13_in,
    input  io_VwirePorts_0_10_13_en,
    output[1:0] io_VwirePorts_0_10_13_out,
    input [1:0] io_VwirePorts_0_10_12_in,
    input  io_VwirePorts_0_10_12_en,
    output[1:0] io_VwirePorts_0_10_12_out,
    input [1:0] io_VwirePorts_0_10_11_in,
    input  io_VwirePorts_0_10_11_en,
    output[1:0] io_VwirePorts_0_10_11_out,
    input [1:0] io_VwirePorts_0_10_10_in,
    input  io_VwirePorts_0_10_10_en,
    output[1:0] io_VwirePorts_0_10_10_out,
    input [1:0] io_VwirePorts_0_10_9_in,
    input  io_VwirePorts_0_10_9_en,
    output[1:0] io_VwirePorts_0_10_9_out,
    input [1:0] io_VwirePorts_0_10_8_in,
    input  io_VwirePorts_0_10_8_en,
    output[1:0] io_VwirePorts_0_10_8_out,
    input [1:0] io_VwirePorts_0_10_7_in,
    input  io_VwirePorts_0_10_7_en,
    output[1:0] io_VwirePorts_0_10_7_out,
    input [1:0] io_VwirePorts_0_10_6_in,
    input  io_VwirePorts_0_10_6_en,
    output[1:0] io_VwirePorts_0_10_6_out,
    input [1:0] io_VwirePorts_0_10_5_in,
    input  io_VwirePorts_0_10_5_en,
    output[1:0] io_VwirePorts_0_10_5_out,
    input [1:0] io_VwirePorts_0_10_4_in,
    input  io_VwirePorts_0_10_4_en,
    output[1:0] io_VwirePorts_0_10_4_out,
    input [1:0] io_VwirePorts_0_10_3_in,
    input  io_VwirePorts_0_10_3_en,
    output[1:0] io_VwirePorts_0_10_3_out,
    input [1:0] io_VwirePorts_0_10_2_in,
    input  io_VwirePorts_0_10_2_en,
    output[1:0] io_VwirePorts_0_10_2_out,
    input [1:0] io_VwirePorts_0_10_1_in,
    input  io_VwirePorts_0_10_1_en,
    output[1:0] io_VwirePorts_0_10_1_out,
    input [1:0] io_VwirePorts_0_10_0_in,
    input  io_VwirePorts_0_10_0_en,
    output[1:0] io_VwirePorts_0_10_0_out,
    input [1:0] io_VwirePorts_0_9_15_in,
    input  io_VwirePorts_0_9_15_en,
    output[1:0] io_VwirePorts_0_9_15_out,
    input [1:0] io_VwirePorts_0_9_14_in,
    input  io_VwirePorts_0_9_14_en,
    output[1:0] io_VwirePorts_0_9_14_out,
    input [1:0] io_VwirePorts_0_9_13_in,
    input  io_VwirePorts_0_9_13_en,
    output[1:0] io_VwirePorts_0_9_13_out,
    input [1:0] io_VwirePorts_0_9_12_in,
    input  io_VwirePorts_0_9_12_en,
    output[1:0] io_VwirePorts_0_9_12_out,
    input [1:0] io_VwirePorts_0_9_11_in,
    input  io_VwirePorts_0_9_11_en,
    output[1:0] io_VwirePorts_0_9_11_out,
    input [1:0] io_VwirePorts_0_9_10_in,
    input  io_VwirePorts_0_9_10_en,
    output[1:0] io_VwirePorts_0_9_10_out,
    input [1:0] io_VwirePorts_0_9_9_in,
    input  io_VwirePorts_0_9_9_en,
    output[1:0] io_VwirePorts_0_9_9_out,
    input [1:0] io_VwirePorts_0_9_8_in,
    input  io_VwirePorts_0_9_8_en,
    output[1:0] io_VwirePorts_0_9_8_out,
    input [1:0] io_VwirePorts_0_9_7_in,
    input  io_VwirePorts_0_9_7_en,
    output[1:0] io_VwirePorts_0_9_7_out,
    input [1:0] io_VwirePorts_0_9_6_in,
    input  io_VwirePorts_0_9_6_en,
    output[1:0] io_VwirePorts_0_9_6_out,
    input [1:0] io_VwirePorts_0_9_5_in,
    input  io_VwirePorts_0_9_5_en,
    output[1:0] io_VwirePorts_0_9_5_out,
    input [1:0] io_VwirePorts_0_9_4_in,
    input  io_VwirePorts_0_9_4_en,
    output[1:0] io_VwirePorts_0_9_4_out,
    input [1:0] io_VwirePorts_0_9_3_in,
    input  io_VwirePorts_0_9_3_en,
    output[1:0] io_VwirePorts_0_9_3_out,
    input [1:0] io_VwirePorts_0_9_2_in,
    input  io_VwirePorts_0_9_2_en,
    output[1:0] io_VwirePorts_0_9_2_out,
    input [1:0] io_VwirePorts_0_9_1_in,
    input  io_VwirePorts_0_9_1_en,
    output[1:0] io_VwirePorts_0_9_1_out,
    input [1:0] io_VwirePorts_0_9_0_in,
    input  io_VwirePorts_0_9_0_en,
    output[1:0] io_VwirePorts_0_9_0_out,
    input [1:0] io_VwirePorts_0_8_15_in,
    input  io_VwirePorts_0_8_15_en,
    output[1:0] io_VwirePorts_0_8_15_out,
    input [1:0] io_VwirePorts_0_8_14_in,
    input  io_VwirePorts_0_8_14_en,
    output[1:0] io_VwirePorts_0_8_14_out,
    input [1:0] io_VwirePorts_0_8_13_in,
    input  io_VwirePorts_0_8_13_en,
    output[1:0] io_VwirePorts_0_8_13_out,
    input [1:0] io_VwirePorts_0_8_12_in,
    input  io_VwirePorts_0_8_12_en,
    output[1:0] io_VwirePorts_0_8_12_out,
    input [1:0] io_VwirePorts_0_8_11_in,
    input  io_VwirePorts_0_8_11_en,
    output[1:0] io_VwirePorts_0_8_11_out,
    input [1:0] io_VwirePorts_0_8_10_in,
    input  io_VwirePorts_0_8_10_en,
    output[1:0] io_VwirePorts_0_8_10_out,
    input [1:0] io_VwirePorts_0_8_9_in,
    input  io_VwirePorts_0_8_9_en,
    output[1:0] io_VwirePorts_0_8_9_out,
    input [1:0] io_VwirePorts_0_8_8_in,
    input  io_VwirePorts_0_8_8_en,
    output[1:0] io_VwirePorts_0_8_8_out,
    input [1:0] io_VwirePorts_0_8_7_in,
    input  io_VwirePorts_0_8_7_en,
    output[1:0] io_VwirePorts_0_8_7_out,
    input [1:0] io_VwirePorts_0_8_6_in,
    input  io_VwirePorts_0_8_6_en,
    output[1:0] io_VwirePorts_0_8_6_out,
    input [1:0] io_VwirePorts_0_8_5_in,
    input  io_VwirePorts_0_8_5_en,
    output[1:0] io_VwirePorts_0_8_5_out,
    input [1:0] io_VwirePorts_0_8_4_in,
    input  io_VwirePorts_0_8_4_en,
    output[1:0] io_VwirePorts_0_8_4_out,
    input [1:0] io_VwirePorts_0_8_3_in,
    input  io_VwirePorts_0_8_3_en,
    output[1:0] io_VwirePorts_0_8_3_out,
    input [1:0] io_VwirePorts_0_8_2_in,
    input  io_VwirePorts_0_8_2_en,
    output[1:0] io_VwirePorts_0_8_2_out,
    input [1:0] io_VwirePorts_0_8_1_in,
    input  io_VwirePorts_0_8_1_en,
    output[1:0] io_VwirePorts_0_8_1_out,
    input [1:0] io_VwirePorts_0_8_0_in,
    input  io_VwirePorts_0_8_0_en,
    output[1:0] io_VwirePorts_0_8_0_out,
    input [1:0] io_VwirePorts_0_7_15_in,
    input  io_VwirePorts_0_7_15_en,
    output[1:0] io_VwirePorts_0_7_15_out,
    input [1:0] io_VwirePorts_0_7_14_in,
    input  io_VwirePorts_0_7_14_en,
    output[1:0] io_VwirePorts_0_7_14_out,
    input [1:0] io_VwirePorts_0_7_13_in,
    input  io_VwirePorts_0_7_13_en,
    output[1:0] io_VwirePorts_0_7_13_out,
    input [1:0] io_VwirePorts_0_7_12_in,
    input  io_VwirePorts_0_7_12_en,
    output[1:0] io_VwirePorts_0_7_12_out,
    input [1:0] io_VwirePorts_0_7_11_in,
    input  io_VwirePorts_0_7_11_en,
    output[1:0] io_VwirePorts_0_7_11_out,
    input [1:0] io_VwirePorts_0_7_10_in,
    input  io_VwirePorts_0_7_10_en,
    output[1:0] io_VwirePorts_0_7_10_out,
    input [1:0] io_VwirePorts_0_7_9_in,
    input  io_VwirePorts_0_7_9_en,
    output[1:0] io_VwirePorts_0_7_9_out,
    input [1:0] io_VwirePorts_0_7_8_in,
    input  io_VwirePorts_0_7_8_en,
    output[1:0] io_VwirePorts_0_7_8_out,
    input [1:0] io_VwirePorts_0_7_7_in,
    input  io_VwirePorts_0_7_7_en,
    output[1:0] io_VwirePorts_0_7_7_out,
    input [1:0] io_VwirePorts_0_7_6_in,
    input  io_VwirePorts_0_7_6_en,
    output[1:0] io_VwirePorts_0_7_6_out,
    input [1:0] io_VwirePorts_0_7_5_in,
    input  io_VwirePorts_0_7_5_en,
    output[1:0] io_VwirePorts_0_7_5_out,
    input [1:0] io_VwirePorts_0_7_4_in,
    input  io_VwirePorts_0_7_4_en,
    output[1:0] io_VwirePorts_0_7_4_out,
    input [1:0] io_VwirePorts_0_7_3_in,
    input  io_VwirePorts_0_7_3_en,
    output[1:0] io_VwirePorts_0_7_3_out,
    input [1:0] io_VwirePorts_0_7_2_in,
    input  io_VwirePorts_0_7_2_en,
    output[1:0] io_VwirePorts_0_7_2_out,
    input [1:0] io_VwirePorts_0_7_1_in,
    input  io_VwirePorts_0_7_1_en,
    output[1:0] io_VwirePorts_0_7_1_out,
    input [1:0] io_VwirePorts_0_7_0_in,
    input  io_VwirePorts_0_7_0_en,
    output[1:0] io_VwirePorts_0_7_0_out,
    input [1:0] io_VwirePorts_0_6_15_in,
    input  io_VwirePorts_0_6_15_en,
    output[1:0] io_VwirePorts_0_6_15_out,
    input [1:0] io_VwirePorts_0_6_14_in,
    input  io_VwirePorts_0_6_14_en,
    output[1:0] io_VwirePorts_0_6_14_out,
    input [1:0] io_VwirePorts_0_6_13_in,
    input  io_VwirePorts_0_6_13_en,
    output[1:0] io_VwirePorts_0_6_13_out,
    input [1:0] io_VwirePorts_0_6_12_in,
    input  io_VwirePorts_0_6_12_en,
    output[1:0] io_VwirePorts_0_6_12_out,
    input [1:0] io_VwirePorts_0_6_11_in,
    input  io_VwirePorts_0_6_11_en,
    output[1:0] io_VwirePorts_0_6_11_out,
    input [1:0] io_VwirePorts_0_6_10_in,
    input  io_VwirePorts_0_6_10_en,
    output[1:0] io_VwirePorts_0_6_10_out,
    input [1:0] io_VwirePorts_0_6_9_in,
    input  io_VwirePorts_0_6_9_en,
    output[1:0] io_VwirePorts_0_6_9_out,
    input [1:0] io_VwirePorts_0_6_8_in,
    input  io_VwirePorts_0_6_8_en,
    output[1:0] io_VwirePorts_0_6_8_out,
    input [1:0] io_VwirePorts_0_6_7_in,
    input  io_VwirePorts_0_6_7_en,
    output[1:0] io_VwirePorts_0_6_7_out,
    input [1:0] io_VwirePorts_0_6_6_in,
    input  io_VwirePorts_0_6_6_en,
    output[1:0] io_VwirePorts_0_6_6_out,
    input [1:0] io_VwirePorts_0_6_5_in,
    input  io_VwirePorts_0_6_5_en,
    output[1:0] io_VwirePorts_0_6_5_out,
    input [1:0] io_VwirePorts_0_6_4_in,
    input  io_VwirePorts_0_6_4_en,
    output[1:0] io_VwirePorts_0_6_4_out,
    input [1:0] io_VwirePorts_0_6_3_in,
    input  io_VwirePorts_0_6_3_en,
    output[1:0] io_VwirePorts_0_6_3_out,
    input [1:0] io_VwirePorts_0_6_2_in,
    input  io_VwirePorts_0_6_2_en,
    output[1:0] io_VwirePorts_0_6_2_out,
    input [1:0] io_VwirePorts_0_6_1_in,
    input  io_VwirePorts_0_6_1_en,
    output[1:0] io_VwirePorts_0_6_1_out,
    input [1:0] io_VwirePorts_0_6_0_in,
    input  io_VwirePorts_0_6_0_en,
    output[1:0] io_VwirePorts_0_6_0_out,
    input [1:0] io_VwirePorts_0_5_15_in,
    input  io_VwirePorts_0_5_15_en,
    output[1:0] io_VwirePorts_0_5_15_out,
    input [1:0] io_VwirePorts_0_5_14_in,
    input  io_VwirePorts_0_5_14_en,
    output[1:0] io_VwirePorts_0_5_14_out,
    input [1:0] io_VwirePorts_0_5_13_in,
    input  io_VwirePorts_0_5_13_en,
    output[1:0] io_VwirePorts_0_5_13_out,
    input [1:0] io_VwirePorts_0_5_12_in,
    input  io_VwirePorts_0_5_12_en,
    output[1:0] io_VwirePorts_0_5_12_out,
    input [1:0] io_VwirePorts_0_5_11_in,
    input  io_VwirePorts_0_5_11_en,
    output[1:0] io_VwirePorts_0_5_11_out,
    input [1:0] io_VwirePorts_0_5_10_in,
    input  io_VwirePorts_0_5_10_en,
    output[1:0] io_VwirePorts_0_5_10_out,
    input [1:0] io_VwirePorts_0_5_9_in,
    input  io_VwirePorts_0_5_9_en,
    output[1:0] io_VwirePorts_0_5_9_out,
    input [1:0] io_VwirePorts_0_5_8_in,
    input  io_VwirePorts_0_5_8_en,
    output[1:0] io_VwirePorts_0_5_8_out,
    input [1:0] io_VwirePorts_0_5_7_in,
    input  io_VwirePorts_0_5_7_en,
    output[1:0] io_VwirePorts_0_5_7_out,
    input [1:0] io_VwirePorts_0_5_6_in,
    input  io_VwirePorts_0_5_6_en,
    output[1:0] io_VwirePorts_0_5_6_out,
    input [1:0] io_VwirePorts_0_5_5_in,
    input  io_VwirePorts_0_5_5_en,
    output[1:0] io_VwirePorts_0_5_5_out,
    input [1:0] io_VwirePorts_0_5_4_in,
    input  io_VwirePorts_0_5_4_en,
    output[1:0] io_VwirePorts_0_5_4_out,
    input [1:0] io_VwirePorts_0_5_3_in,
    input  io_VwirePorts_0_5_3_en,
    output[1:0] io_VwirePorts_0_5_3_out,
    input [1:0] io_VwirePorts_0_5_2_in,
    input  io_VwirePorts_0_5_2_en,
    output[1:0] io_VwirePorts_0_5_2_out,
    input [1:0] io_VwirePorts_0_5_1_in,
    input  io_VwirePorts_0_5_1_en,
    output[1:0] io_VwirePorts_0_5_1_out,
    input [1:0] io_VwirePorts_0_5_0_in,
    input  io_VwirePorts_0_5_0_en,
    output[1:0] io_VwirePorts_0_5_0_out,
    input [1:0] io_VwirePorts_0_4_15_in,
    input  io_VwirePorts_0_4_15_en,
    output[1:0] io_VwirePorts_0_4_15_out,
    input [1:0] io_VwirePorts_0_4_14_in,
    input  io_VwirePorts_0_4_14_en,
    output[1:0] io_VwirePorts_0_4_14_out,
    input [1:0] io_VwirePorts_0_4_13_in,
    input  io_VwirePorts_0_4_13_en,
    output[1:0] io_VwirePorts_0_4_13_out,
    input [1:0] io_VwirePorts_0_4_12_in,
    input  io_VwirePorts_0_4_12_en,
    output[1:0] io_VwirePorts_0_4_12_out,
    input [1:0] io_VwirePorts_0_4_11_in,
    input  io_VwirePorts_0_4_11_en,
    output[1:0] io_VwirePorts_0_4_11_out,
    input [1:0] io_VwirePorts_0_4_10_in,
    input  io_VwirePorts_0_4_10_en,
    output[1:0] io_VwirePorts_0_4_10_out,
    input [1:0] io_VwirePorts_0_4_9_in,
    input  io_VwirePorts_0_4_9_en,
    output[1:0] io_VwirePorts_0_4_9_out,
    input [1:0] io_VwirePorts_0_4_8_in,
    input  io_VwirePorts_0_4_8_en,
    output[1:0] io_VwirePorts_0_4_8_out,
    input [1:0] io_VwirePorts_0_4_7_in,
    input  io_VwirePorts_0_4_7_en,
    output[1:0] io_VwirePorts_0_4_7_out,
    input [1:0] io_VwirePorts_0_4_6_in,
    input  io_VwirePorts_0_4_6_en,
    output[1:0] io_VwirePorts_0_4_6_out,
    input [1:0] io_VwirePorts_0_4_5_in,
    input  io_VwirePorts_0_4_5_en,
    output[1:0] io_VwirePorts_0_4_5_out,
    input [1:0] io_VwirePorts_0_4_4_in,
    input  io_VwirePorts_0_4_4_en,
    output[1:0] io_VwirePorts_0_4_4_out,
    input [1:0] io_VwirePorts_0_4_3_in,
    input  io_VwirePorts_0_4_3_en,
    output[1:0] io_VwirePorts_0_4_3_out,
    input [1:0] io_VwirePorts_0_4_2_in,
    input  io_VwirePorts_0_4_2_en,
    output[1:0] io_VwirePorts_0_4_2_out,
    input [1:0] io_VwirePorts_0_4_1_in,
    input  io_VwirePorts_0_4_1_en,
    output[1:0] io_VwirePorts_0_4_1_out,
    input [1:0] io_VwirePorts_0_4_0_in,
    input  io_VwirePorts_0_4_0_en,
    output[1:0] io_VwirePorts_0_4_0_out,
    input [1:0] io_VwirePorts_0_3_15_in,
    input  io_VwirePorts_0_3_15_en,
    output[1:0] io_VwirePorts_0_3_15_out,
    input [1:0] io_VwirePorts_0_3_14_in,
    input  io_VwirePorts_0_3_14_en,
    output[1:0] io_VwirePorts_0_3_14_out,
    input [1:0] io_VwirePorts_0_3_13_in,
    input  io_VwirePorts_0_3_13_en,
    output[1:0] io_VwirePorts_0_3_13_out,
    input [1:0] io_VwirePorts_0_3_12_in,
    input  io_VwirePorts_0_3_12_en,
    output[1:0] io_VwirePorts_0_3_12_out,
    input [1:0] io_VwirePorts_0_3_11_in,
    input  io_VwirePorts_0_3_11_en,
    output[1:0] io_VwirePorts_0_3_11_out,
    input [1:0] io_VwirePorts_0_3_10_in,
    input  io_VwirePorts_0_3_10_en,
    output[1:0] io_VwirePorts_0_3_10_out,
    input [1:0] io_VwirePorts_0_3_9_in,
    input  io_VwirePorts_0_3_9_en,
    output[1:0] io_VwirePorts_0_3_9_out,
    input [1:0] io_VwirePorts_0_3_8_in,
    input  io_VwirePorts_0_3_8_en,
    output[1:0] io_VwirePorts_0_3_8_out,
    input [1:0] io_VwirePorts_0_3_7_in,
    input  io_VwirePorts_0_3_7_en,
    output[1:0] io_VwirePorts_0_3_7_out,
    input [1:0] io_VwirePorts_0_3_6_in,
    input  io_VwirePorts_0_3_6_en,
    output[1:0] io_VwirePorts_0_3_6_out,
    input [1:0] io_VwirePorts_0_3_5_in,
    input  io_VwirePorts_0_3_5_en,
    output[1:0] io_VwirePorts_0_3_5_out,
    input [1:0] io_VwirePorts_0_3_4_in,
    input  io_VwirePorts_0_3_4_en,
    output[1:0] io_VwirePorts_0_3_4_out,
    input [1:0] io_VwirePorts_0_3_3_in,
    input  io_VwirePorts_0_3_3_en,
    output[1:0] io_VwirePorts_0_3_3_out,
    input [1:0] io_VwirePorts_0_3_2_in,
    input  io_VwirePorts_0_3_2_en,
    output[1:0] io_VwirePorts_0_3_2_out,
    input [1:0] io_VwirePorts_0_3_1_in,
    input  io_VwirePorts_0_3_1_en,
    output[1:0] io_VwirePorts_0_3_1_out,
    input [1:0] io_VwirePorts_0_3_0_in,
    input  io_VwirePorts_0_3_0_en,
    output[1:0] io_VwirePorts_0_3_0_out,
    input [1:0] io_VwirePorts_0_2_15_in,
    input  io_VwirePorts_0_2_15_en,
    output[1:0] io_VwirePorts_0_2_15_out,
    input [1:0] io_VwirePorts_0_2_14_in,
    input  io_VwirePorts_0_2_14_en,
    output[1:0] io_VwirePorts_0_2_14_out,
    input [1:0] io_VwirePorts_0_2_13_in,
    input  io_VwirePorts_0_2_13_en,
    output[1:0] io_VwirePorts_0_2_13_out,
    input [1:0] io_VwirePorts_0_2_12_in,
    input  io_VwirePorts_0_2_12_en,
    output[1:0] io_VwirePorts_0_2_12_out,
    input [1:0] io_VwirePorts_0_2_11_in,
    input  io_VwirePorts_0_2_11_en,
    output[1:0] io_VwirePorts_0_2_11_out,
    input [1:0] io_VwirePorts_0_2_10_in,
    input  io_VwirePorts_0_2_10_en,
    output[1:0] io_VwirePorts_0_2_10_out,
    input [1:0] io_VwirePorts_0_2_9_in,
    input  io_VwirePorts_0_2_9_en,
    output[1:0] io_VwirePorts_0_2_9_out,
    input [1:0] io_VwirePorts_0_2_8_in,
    input  io_VwirePorts_0_2_8_en,
    output[1:0] io_VwirePorts_0_2_8_out,
    input [1:0] io_VwirePorts_0_2_7_in,
    input  io_VwirePorts_0_2_7_en,
    output[1:0] io_VwirePorts_0_2_7_out,
    input [1:0] io_VwirePorts_0_2_6_in,
    input  io_VwirePorts_0_2_6_en,
    output[1:0] io_VwirePorts_0_2_6_out,
    input [1:0] io_VwirePorts_0_2_5_in,
    input  io_VwirePorts_0_2_5_en,
    output[1:0] io_VwirePorts_0_2_5_out,
    input [1:0] io_VwirePorts_0_2_4_in,
    input  io_VwirePorts_0_2_4_en,
    output[1:0] io_VwirePorts_0_2_4_out,
    input [1:0] io_VwirePorts_0_2_3_in,
    input  io_VwirePorts_0_2_3_en,
    output[1:0] io_VwirePorts_0_2_3_out,
    input [1:0] io_VwirePorts_0_2_2_in,
    input  io_VwirePorts_0_2_2_en,
    output[1:0] io_VwirePorts_0_2_2_out,
    input [1:0] io_VwirePorts_0_2_1_in,
    input  io_VwirePorts_0_2_1_en,
    output[1:0] io_VwirePorts_0_2_1_out,
    input [1:0] io_VwirePorts_0_2_0_in,
    input  io_VwirePorts_0_2_0_en,
    output[1:0] io_VwirePorts_0_2_0_out,
    input [1:0] io_VwirePorts_0_1_15_in,
    input  io_VwirePorts_0_1_15_en,
    output[1:0] io_VwirePorts_0_1_15_out,
    input [1:0] io_VwirePorts_0_1_14_in,
    input  io_VwirePorts_0_1_14_en,
    output[1:0] io_VwirePorts_0_1_14_out,
    input [1:0] io_VwirePorts_0_1_13_in,
    input  io_VwirePorts_0_1_13_en,
    output[1:0] io_VwirePorts_0_1_13_out,
    input [1:0] io_VwirePorts_0_1_12_in,
    input  io_VwirePorts_0_1_12_en,
    output[1:0] io_VwirePorts_0_1_12_out,
    input [1:0] io_VwirePorts_0_1_11_in,
    input  io_VwirePorts_0_1_11_en,
    output[1:0] io_VwirePorts_0_1_11_out,
    input [1:0] io_VwirePorts_0_1_10_in,
    input  io_VwirePorts_0_1_10_en,
    output[1:0] io_VwirePorts_0_1_10_out,
    input [1:0] io_VwirePorts_0_1_9_in,
    input  io_VwirePorts_0_1_9_en,
    output[1:0] io_VwirePorts_0_1_9_out,
    input [1:0] io_VwirePorts_0_1_8_in,
    input  io_VwirePorts_0_1_8_en,
    output[1:0] io_VwirePorts_0_1_8_out,
    input [1:0] io_VwirePorts_0_1_7_in,
    input  io_VwirePorts_0_1_7_en,
    output[1:0] io_VwirePorts_0_1_7_out,
    input [1:0] io_VwirePorts_0_1_6_in,
    input  io_VwirePorts_0_1_6_en,
    output[1:0] io_VwirePorts_0_1_6_out,
    input [1:0] io_VwirePorts_0_1_5_in,
    input  io_VwirePorts_0_1_5_en,
    output[1:0] io_VwirePorts_0_1_5_out,
    input [1:0] io_VwirePorts_0_1_4_in,
    input  io_VwirePorts_0_1_4_en,
    output[1:0] io_VwirePorts_0_1_4_out,
    input [1:0] io_VwirePorts_0_1_3_in,
    input  io_VwirePorts_0_1_3_en,
    output[1:0] io_VwirePorts_0_1_3_out,
    input [1:0] io_VwirePorts_0_1_2_in,
    input  io_VwirePorts_0_1_2_en,
    output[1:0] io_VwirePorts_0_1_2_out,
    input [1:0] io_VwirePorts_0_1_1_in,
    input  io_VwirePorts_0_1_1_en,
    output[1:0] io_VwirePorts_0_1_1_out,
    input [1:0] io_VwirePorts_0_1_0_in,
    input  io_VwirePorts_0_1_0_en,
    output[1:0] io_VwirePorts_0_1_0_out,
    input [1:0] io_VwirePorts_0_0_15_in,
    input  io_VwirePorts_0_0_15_en,
    output[1:0] io_VwirePorts_0_0_15_out,
    input [1:0] io_VwirePorts_0_0_14_in,
    input  io_VwirePorts_0_0_14_en,
    output[1:0] io_VwirePorts_0_0_14_out,
    input [1:0] io_VwirePorts_0_0_13_in,
    input  io_VwirePorts_0_0_13_en,
    output[1:0] io_VwirePorts_0_0_13_out,
    input [1:0] io_VwirePorts_0_0_12_in,
    input  io_VwirePorts_0_0_12_en,
    output[1:0] io_VwirePorts_0_0_12_out,
    input [1:0] io_VwirePorts_0_0_11_in,
    input  io_VwirePorts_0_0_11_en,
    output[1:0] io_VwirePorts_0_0_11_out,
    input [1:0] io_VwirePorts_0_0_10_in,
    input  io_VwirePorts_0_0_10_en,
    output[1:0] io_VwirePorts_0_0_10_out,
    input [1:0] io_VwirePorts_0_0_9_in,
    input  io_VwirePorts_0_0_9_en,
    output[1:0] io_VwirePorts_0_0_9_out,
    input [1:0] io_VwirePorts_0_0_8_in,
    input  io_VwirePorts_0_0_8_en,
    output[1:0] io_VwirePorts_0_0_8_out,
    input [1:0] io_VwirePorts_0_0_7_in,
    input  io_VwirePorts_0_0_7_en,
    output[1:0] io_VwirePorts_0_0_7_out,
    input [1:0] io_VwirePorts_0_0_6_in,
    input  io_VwirePorts_0_0_6_en,
    output[1:0] io_VwirePorts_0_0_6_out,
    input [1:0] io_VwirePorts_0_0_5_in,
    input  io_VwirePorts_0_0_5_en,
    output[1:0] io_VwirePorts_0_0_5_out,
    input [1:0] io_VwirePorts_0_0_4_in,
    input  io_VwirePorts_0_0_4_en,
    output[1:0] io_VwirePorts_0_0_4_out,
    input [1:0] io_VwirePorts_0_0_3_in,
    input  io_VwirePorts_0_0_3_en,
    output[1:0] io_VwirePorts_0_0_3_out,
    input [1:0] io_VwirePorts_0_0_2_in,
    input  io_VwirePorts_0_0_2_en,
    output[1:0] io_VwirePorts_0_0_2_out,
    input [1:0] io_VwirePorts_0_0_1_in,
    input  io_VwirePorts_0_0_1_en,
    output[1:0] io_VwirePorts_0_0_1_out,
    input [1:0] io_VwirePorts_0_0_0_in,
    input  io_VwirePorts_0_0_0_en,
    output[1:0] io_VwirePorts_0_0_0_out
);

  wire[1:0] Vwire_io_out;
  wire[1:0] Vwire_1_io_out;
  wire[1:0] Vwire_2_io_out;
  wire[1:0] Vwire_3_io_out;
  wire[1:0] Vwire_4_io_out;
  wire[1:0] Vwire_5_io_out;
  wire[1:0] Vwire_6_io_out;
  wire[1:0] Vwire_7_io_out;
  wire[1:0] Vwire_8_io_out;
  wire[1:0] Vwire_9_io_out;
  wire[1:0] Vwire_10_io_out;
  wire[1:0] Vwire_11_io_out;
  wire[1:0] Vwire_12_io_out;
  wire[1:0] Vwire_13_io_out;
  wire[1:0] Vwire_14_io_out;
  wire[1:0] Vwire_15_io_out;
  wire[1:0] Vwire_16_io_out;
  wire[1:0] Vwire_17_io_out;
  wire[1:0] Vwire_18_io_out;
  wire[1:0] Vwire_19_io_out;
  wire[1:0] Vwire_20_io_out;
  wire[1:0] Vwire_21_io_out;
  wire[1:0] Vwire_22_io_out;
  wire[1:0] Vwire_23_io_out;
  wire[1:0] Vwire_24_io_out;
  wire[1:0] Vwire_25_io_out;
  wire[1:0] Vwire_26_io_out;
  wire[1:0] Vwire_27_io_out;
  wire[1:0] Vwire_28_io_out;
  wire[1:0] Vwire_29_io_out;
  wire[1:0] Vwire_30_io_out;
  wire[1:0] Vwire_31_io_out;
  wire[1:0] Vwire_32_io_out;
  wire[1:0] Vwire_33_io_out;
  wire[1:0] Vwire_34_io_out;
  wire[1:0] Vwire_35_io_out;
  wire[1:0] Vwire_36_io_out;
  wire[1:0] Vwire_37_io_out;
  wire[1:0] Vwire_38_io_out;
  wire[1:0] Vwire_39_io_out;
  wire[1:0] Vwire_40_io_out;
  wire[1:0] Vwire_41_io_out;
  wire[1:0] Vwire_42_io_out;
  wire[1:0] Vwire_43_io_out;
  wire[1:0] Vwire_44_io_out;
  wire[1:0] Vwire_45_io_out;
  wire[1:0] Vwire_46_io_out;
  wire[1:0] Vwire_47_io_out;
  wire[1:0] Vwire_48_io_out;
  wire[1:0] Vwire_49_io_out;
  wire[1:0] Vwire_50_io_out;
  wire[1:0] Vwire_51_io_out;
  wire[1:0] Vwire_52_io_out;
  wire[1:0] Vwire_53_io_out;
  wire[1:0] Vwire_54_io_out;
  wire[1:0] Vwire_55_io_out;
  wire[1:0] Vwire_56_io_out;
  wire[1:0] Vwire_57_io_out;
  wire[1:0] Vwire_58_io_out;
  wire[1:0] Vwire_59_io_out;
  wire[1:0] Vwire_60_io_out;
  wire[1:0] Vwire_61_io_out;
  wire[1:0] Vwire_62_io_out;
  wire[1:0] Vwire_63_io_out;
  wire[1:0] Vwire_64_io_out;
  wire[1:0] Vwire_65_io_out;
  wire[1:0] Vwire_66_io_out;
  wire[1:0] Vwire_67_io_out;
  wire[1:0] Vwire_68_io_out;
  wire[1:0] Vwire_69_io_out;
  wire[1:0] Vwire_70_io_out;
  wire[1:0] Vwire_71_io_out;
  wire[1:0] Vwire_72_io_out;
  wire[1:0] Vwire_73_io_out;
  wire[1:0] Vwire_74_io_out;
  wire[1:0] Vwire_75_io_out;
  wire[1:0] Vwire_76_io_out;
  wire[1:0] Vwire_77_io_out;
  wire[1:0] Vwire_78_io_out;
  wire[1:0] Vwire_79_io_out;
  wire[1:0] Vwire_80_io_out;
  wire[1:0] Vwire_81_io_out;
  wire[1:0] Vwire_82_io_out;
  wire[1:0] Vwire_83_io_out;
  wire[1:0] Vwire_84_io_out;
  wire[1:0] Vwire_85_io_out;
  wire[1:0] Vwire_86_io_out;
  wire[1:0] Vwire_87_io_out;
  wire[1:0] Vwire_88_io_out;
  wire[1:0] Vwire_89_io_out;
  wire[1:0] Vwire_90_io_out;
  wire[1:0] Vwire_91_io_out;
  wire[1:0] Vwire_92_io_out;
  wire[1:0] Vwire_93_io_out;
  wire[1:0] Vwire_94_io_out;
  wire[1:0] Vwire_95_io_out;
  wire[1:0] Vwire_96_io_out;
  wire[1:0] Vwire_97_io_out;
  wire[1:0] Vwire_98_io_out;
  wire[1:0] Vwire_99_io_out;
  wire[1:0] Vwire_100_io_out;
  wire[1:0] Vwire_101_io_out;
  wire[1:0] Vwire_102_io_out;
  wire[1:0] Vwire_103_io_out;
  wire[1:0] Vwire_104_io_out;
  wire[1:0] Vwire_105_io_out;
  wire[1:0] Vwire_106_io_out;
  wire[1:0] Vwire_107_io_out;
  wire[1:0] Vwire_108_io_out;
  wire[1:0] Vwire_109_io_out;
  wire[1:0] Vwire_110_io_out;
  wire[1:0] Vwire_111_io_out;
  wire[1:0] Vwire_112_io_out;
  wire[1:0] Vwire_113_io_out;
  wire[1:0] Vwire_114_io_out;
  wire[1:0] Vwire_115_io_out;
  wire[1:0] Vwire_116_io_out;
  wire[1:0] Vwire_117_io_out;
  wire[1:0] Vwire_118_io_out;
  wire[1:0] Vwire_119_io_out;
  wire[1:0] Vwire_120_io_out;
  wire[1:0] Vwire_121_io_out;
  wire[1:0] Vwire_122_io_out;
  wire[1:0] Vwire_123_io_out;
  wire[1:0] Vwire_124_io_out;
  wire[1:0] Vwire_125_io_out;
  wire[1:0] Vwire_126_io_out;
  wire[1:0] Vwire_127_io_out;
  wire[1:0] Vwire_128_io_out;
  wire[1:0] Vwire_129_io_out;
  wire[1:0] Vwire_130_io_out;
  wire[1:0] Vwire_131_io_out;
  wire[1:0] Vwire_132_io_out;
  wire[1:0] Vwire_133_io_out;
  wire[1:0] Vwire_134_io_out;
  wire[1:0] Vwire_135_io_out;
  wire[1:0] Vwire_136_io_out;
  wire[1:0] Vwire_137_io_out;
  wire[1:0] Vwire_138_io_out;
  wire[1:0] Vwire_139_io_out;
  wire[1:0] Vwire_140_io_out;
  wire[1:0] Vwire_141_io_out;
  wire[1:0] Vwire_142_io_out;
  wire[1:0] Vwire_143_io_out;
  wire[1:0] Vwire_144_io_out;
  wire[1:0] Vwire_145_io_out;
  wire[1:0] Vwire_146_io_out;
  wire[1:0] Vwire_147_io_out;
  wire[1:0] Vwire_148_io_out;
  wire[1:0] Vwire_149_io_out;
  wire[1:0] Vwire_150_io_out;
  wire[1:0] Vwire_151_io_out;
  wire[1:0] Vwire_152_io_out;
  wire[1:0] Vwire_153_io_out;
  wire[1:0] Vwire_154_io_out;
  wire[1:0] Vwire_155_io_out;
  wire[1:0] Vwire_156_io_out;
  wire[1:0] Vwire_157_io_out;
  wire[1:0] Vwire_158_io_out;
  wire[1:0] Vwire_159_io_out;
  wire[1:0] Vwire_160_io_out;
  wire[1:0] Vwire_161_io_out;
  wire[1:0] Vwire_162_io_out;
  wire[1:0] Vwire_163_io_out;
  wire[1:0] Vwire_164_io_out;
  wire[1:0] Vwire_165_io_out;
  wire[1:0] Vwire_166_io_out;
  wire[1:0] Vwire_167_io_out;
  wire[1:0] Vwire_168_io_out;
  wire[1:0] Vwire_169_io_out;
  wire[1:0] Vwire_170_io_out;
  wire[1:0] Vwire_171_io_out;
  wire[1:0] Vwire_172_io_out;
  wire[1:0] Vwire_173_io_out;
  wire[1:0] Vwire_174_io_out;
  wire[1:0] Vwire_175_io_out;
  wire[1:0] Vwire_176_io_out;
  wire[1:0] Vwire_177_io_out;
  wire[1:0] Vwire_178_io_out;
  wire[1:0] Vwire_179_io_out;
  wire[1:0] Vwire_180_io_out;
  wire[1:0] Vwire_181_io_out;
  wire[1:0] Vwire_182_io_out;
  wire[1:0] Vwire_183_io_out;


`ifndef SYNTHESIS
// synthesis translate_off
  assign io_VwirePorts_0_0_2_out = {1{$random}};
  assign io_VwirePorts_0_0_6_out = {1{$random}};
  assign io_VwirePorts_0_0_7_out = {1{$random}};
  assign io_VwirePorts_0_0_8_out = {1{$random}};
  assign io_VwirePorts_0_0_9_out = {1{$random}};
  assign io_VwirePorts_0_0_10_out = {1{$random}};
  assign io_VwirePorts_0_0_11_out = {1{$random}};
  assign io_VwirePorts_0_0_12_out = {1{$random}};
  assign io_VwirePorts_0_0_13_out = {1{$random}};
  assign io_VwirePorts_0_0_14_out = {1{$random}};
  assign io_VwirePorts_0_0_15_out = {1{$random}};
  assign io_VwirePorts_0_1_2_out = {1{$random}};
  assign io_VwirePorts_0_1_6_out = {1{$random}};
  assign io_VwirePorts_0_1_7_out = {1{$random}};
  assign io_VwirePorts_0_1_8_out = {1{$random}};
  assign io_VwirePorts_0_1_9_out = {1{$random}};
  assign io_VwirePorts_0_1_10_out = {1{$random}};
  assign io_VwirePorts_0_1_11_out = {1{$random}};
  assign io_VwirePorts_0_1_12_out = {1{$random}};
  assign io_VwirePorts_0_1_13_out = {1{$random}};
  assign io_VwirePorts_0_1_14_out = {1{$random}};
  assign io_VwirePorts_0_1_15_out = {1{$random}};
  assign io_VwirePorts_0_2_2_out = {1{$random}};
  assign io_VwirePorts_0_2_6_out = {1{$random}};
  assign io_VwirePorts_0_2_7_out = {1{$random}};
  assign io_VwirePorts_0_2_8_out = {1{$random}};
  assign io_VwirePorts_0_2_9_out = {1{$random}};
  assign io_VwirePorts_0_2_10_out = {1{$random}};
  assign io_VwirePorts_0_2_11_out = {1{$random}};
  assign io_VwirePorts_0_2_12_out = {1{$random}};
  assign io_VwirePorts_0_2_13_out = {1{$random}};
  assign io_VwirePorts_0_2_14_out = {1{$random}};
  assign io_VwirePorts_0_2_15_out = {1{$random}};
  assign io_VwirePorts_0_3_2_out = {1{$random}};
  assign io_VwirePorts_0_3_6_out = {1{$random}};
  assign io_VwirePorts_0_3_7_out = {1{$random}};
  assign io_VwirePorts_0_3_8_out = {1{$random}};
  assign io_VwirePorts_0_3_9_out = {1{$random}};
  assign io_VwirePorts_0_3_10_out = {1{$random}};
  assign io_VwirePorts_0_3_11_out = {1{$random}};
  assign io_VwirePorts_0_3_12_out = {1{$random}};
  assign io_VwirePorts_0_3_13_out = {1{$random}};
  assign io_VwirePorts_0_3_14_out = {1{$random}};
  assign io_VwirePorts_0_3_15_out = {1{$random}};
  assign io_VwirePorts_0_4_2_out = {1{$random}};
  assign io_VwirePorts_0_4_6_out = {1{$random}};
  assign io_VwirePorts_0_4_7_out = {1{$random}};
  assign io_VwirePorts_0_4_8_out = {1{$random}};
  assign io_VwirePorts_0_4_9_out = {1{$random}};
  assign io_VwirePorts_0_4_10_out = {1{$random}};
  assign io_VwirePorts_0_4_11_out = {1{$random}};
  assign io_VwirePorts_0_4_12_out = {1{$random}};
  assign io_VwirePorts_0_4_13_out = {1{$random}};
  assign io_VwirePorts_0_4_14_out = {1{$random}};
  assign io_VwirePorts_0_4_15_out = {1{$random}};
  assign io_VwirePorts_0_5_2_out = {1{$random}};
  assign io_VwirePorts_0_5_6_out = {1{$random}};
  assign io_VwirePorts_0_5_7_out = {1{$random}};
  assign io_VwirePorts_0_5_8_out = {1{$random}};
  assign io_VwirePorts_0_5_9_out = {1{$random}};
  assign io_VwirePorts_0_5_10_out = {1{$random}};
  assign io_VwirePorts_0_5_11_out = {1{$random}};
  assign io_VwirePorts_0_5_12_out = {1{$random}};
  assign io_VwirePorts_0_5_13_out = {1{$random}};
  assign io_VwirePorts_0_5_14_out = {1{$random}};
  assign io_VwirePorts_0_5_15_out = {1{$random}};
  assign io_VwirePorts_0_6_2_out = {1{$random}};
  assign io_VwirePorts_0_6_6_out = {1{$random}};
  assign io_VwirePorts_0_6_7_out = {1{$random}};
  assign io_VwirePorts_0_6_8_out = {1{$random}};
  assign io_VwirePorts_0_6_9_out = {1{$random}};
  assign io_VwirePorts_0_6_10_out = {1{$random}};
  assign io_VwirePorts_0_6_11_out = {1{$random}};
  assign io_VwirePorts_0_6_12_out = {1{$random}};
  assign io_VwirePorts_0_6_13_out = {1{$random}};
  assign io_VwirePorts_0_6_14_out = {1{$random}};
  assign io_VwirePorts_0_6_15_out = {1{$random}};
  assign io_VwirePorts_0_7_2_out = {1{$random}};
  assign io_VwirePorts_0_7_6_out = {1{$random}};
  assign io_VwirePorts_0_7_7_out = {1{$random}};
  assign io_VwirePorts_0_7_8_out = {1{$random}};
  assign io_VwirePorts_0_7_9_out = {1{$random}};
  assign io_VwirePorts_0_7_10_out = {1{$random}};
  assign io_VwirePorts_0_7_11_out = {1{$random}};
  assign io_VwirePorts_0_7_12_out = {1{$random}};
  assign io_VwirePorts_0_7_13_out = {1{$random}};
  assign io_VwirePorts_0_7_14_out = {1{$random}};
  assign io_VwirePorts_0_7_15_out = {1{$random}};
  assign io_VwirePorts_0_8_2_out = {1{$random}};
  assign io_VwirePorts_0_8_6_out = {1{$random}};
  assign io_VwirePorts_0_8_7_out = {1{$random}};
  assign io_VwirePorts_0_8_8_out = {1{$random}};
  assign io_VwirePorts_0_8_9_out = {1{$random}};
  assign io_VwirePorts_0_8_10_out = {1{$random}};
  assign io_VwirePorts_0_8_11_out = {1{$random}};
  assign io_VwirePorts_0_8_12_out = {1{$random}};
  assign io_VwirePorts_0_8_13_out = {1{$random}};
  assign io_VwirePorts_0_8_14_out = {1{$random}};
  assign io_VwirePorts_0_8_15_out = {1{$random}};
  assign io_VwirePorts_0_9_2_out = {1{$random}};
  assign io_VwirePorts_0_9_6_out = {1{$random}};
  assign io_VwirePorts_0_9_7_out = {1{$random}};
  assign io_VwirePorts_0_9_8_out = {1{$random}};
  assign io_VwirePorts_0_9_9_out = {1{$random}};
  assign io_VwirePorts_0_9_10_out = {1{$random}};
  assign io_VwirePorts_0_9_11_out = {1{$random}};
  assign io_VwirePorts_0_9_12_out = {1{$random}};
  assign io_VwirePorts_0_9_13_out = {1{$random}};
  assign io_VwirePorts_0_9_14_out = {1{$random}};
  assign io_VwirePorts_0_9_15_out = {1{$random}};
  assign io_VwirePorts_0_10_2_out = {1{$random}};
  assign io_VwirePorts_0_10_6_out = {1{$random}};
  assign io_VwirePorts_0_10_7_out = {1{$random}};
  assign io_VwirePorts_0_10_8_out = {1{$random}};
  assign io_VwirePorts_0_10_9_out = {1{$random}};
  assign io_VwirePorts_0_10_10_out = {1{$random}};
  assign io_VwirePorts_0_10_11_out = {1{$random}};
  assign io_VwirePorts_0_10_12_out = {1{$random}};
  assign io_VwirePorts_0_10_13_out = {1{$random}};
  assign io_VwirePorts_0_10_14_out = {1{$random}};
  assign io_VwirePorts_0_10_15_out = {1{$random}};
  assign io_VwirePorts_0_11_2_out = {1{$random}};
  assign io_VwirePorts_0_11_6_out = {1{$random}};
  assign io_VwirePorts_0_11_7_out = {1{$random}};
  assign io_VwirePorts_0_11_8_out = {1{$random}};
  assign io_VwirePorts_0_11_9_out = {1{$random}};
  assign io_VwirePorts_0_11_10_out = {1{$random}};
  assign io_VwirePorts_0_11_11_out = {1{$random}};
  assign io_VwirePorts_0_11_12_out = {1{$random}};
  assign io_VwirePorts_0_11_13_out = {1{$random}};
  assign io_VwirePorts_0_11_14_out = {1{$random}};
  assign io_VwirePorts_0_11_15_out = {1{$random}};
  assign io_VwirePorts_0_12_2_out = {1{$random}};
  assign io_VwirePorts_0_12_6_out = {1{$random}};
  assign io_VwirePorts_0_12_7_out = {1{$random}};
  assign io_VwirePorts_0_12_8_out = {1{$random}};
  assign io_VwirePorts_0_12_9_out = {1{$random}};
  assign io_VwirePorts_0_12_10_out = {1{$random}};
  assign io_VwirePorts_0_12_11_out = {1{$random}};
  assign io_VwirePorts_0_12_12_out = {1{$random}};
  assign io_VwirePorts_0_12_13_out = {1{$random}};
  assign io_VwirePorts_0_12_14_out = {1{$random}};
  assign io_VwirePorts_0_12_15_out = {1{$random}};
  assign io_VwirePorts_0_13_2_out = {1{$random}};
  assign io_VwirePorts_0_13_6_out = {1{$random}};
  assign io_VwirePorts_0_13_7_out = {1{$random}};
  assign io_VwirePorts_0_13_8_out = {1{$random}};
  assign io_VwirePorts_0_13_9_out = {1{$random}};
  assign io_VwirePorts_0_13_10_out = {1{$random}};
  assign io_VwirePorts_0_13_11_out = {1{$random}};
  assign io_VwirePorts_0_13_12_out = {1{$random}};
  assign io_VwirePorts_0_13_13_out = {1{$random}};
  assign io_VwirePorts_0_13_14_out = {1{$random}};
  assign io_VwirePorts_0_13_15_out = {1{$random}};
  assign io_VwirePorts_0_14_2_out = {1{$random}};
  assign io_VwirePorts_0_14_6_out = {1{$random}};
  assign io_VwirePorts_0_14_7_out = {1{$random}};
  assign io_VwirePorts_0_14_8_out = {1{$random}};
  assign io_VwirePorts_0_14_9_out = {1{$random}};
  assign io_VwirePorts_0_14_10_out = {1{$random}};
  assign io_VwirePorts_0_14_11_out = {1{$random}};
  assign io_VwirePorts_0_14_12_out = {1{$random}};
  assign io_VwirePorts_0_14_13_out = {1{$random}};
  assign io_VwirePorts_0_14_14_out = {1{$random}};
  assign io_VwirePorts_0_14_15_out = {1{$random}};
  assign io_VwirePorts_0_15_2_out = {1{$random}};
  assign io_VwirePorts_0_15_6_out = {1{$random}};
  assign io_VwirePorts_0_15_7_out = {1{$random}};
  assign io_VwirePorts_0_15_8_out = {1{$random}};
  assign io_VwirePorts_0_15_9_out = {1{$random}};
  assign io_VwirePorts_0_15_10_out = {1{$random}};
  assign io_VwirePorts_0_15_11_out = {1{$random}};
  assign io_VwirePorts_0_15_12_out = {1{$random}};
  assign io_VwirePorts_0_15_13_out = {1{$random}};
  assign io_VwirePorts_0_15_14_out = {1{$random}};
  assign io_VwirePorts_0_15_15_out = {1{$random}};
  assign io_VwirePorts_0_16_2_out = {1{$random}};
  assign io_VwirePorts_0_16_6_out = {1{$random}};
  assign io_VwirePorts_0_16_7_out = {1{$random}};
  assign io_VwirePorts_0_16_8_out = {1{$random}};
  assign io_VwirePorts_0_16_9_out = {1{$random}};
  assign io_VwirePorts_0_16_10_out = {1{$random}};
  assign io_VwirePorts_0_16_11_out = {1{$random}};
  assign io_VwirePorts_0_16_12_out = {1{$random}};
  assign io_VwirePorts_0_16_13_out = {1{$random}};
  assign io_VwirePorts_0_16_14_out = {1{$random}};
  assign io_VwirePorts_0_16_15_out = {1{$random}};
  assign io_VwirePorts_0_17_2_out = {1{$random}};
  assign io_VwirePorts_0_17_6_out = {1{$random}};
  assign io_VwirePorts_0_17_7_out = {1{$random}};
  assign io_VwirePorts_0_17_8_out = {1{$random}};
  assign io_VwirePorts_0_17_9_out = {1{$random}};
  assign io_VwirePorts_0_17_10_out = {1{$random}};
  assign io_VwirePorts_0_17_11_out = {1{$random}};
  assign io_VwirePorts_0_17_12_out = {1{$random}};
  assign io_VwirePorts_0_17_13_out = {1{$random}};
  assign io_VwirePorts_0_17_14_out = {1{$random}};
  assign io_VwirePorts_0_17_15_out = {1{$random}};
  assign io_VwirePorts_0_18_2_out = {1{$random}};
  assign io_VwirePorts_0_18_6_out = {1{$random}};
  assign io_VwirePorts_0_18_7_out = {1{$random}};
  assign io_VwirePorts_0_18_8_out = {1{$random}};
  assign io_VwirePorts_0_18_9_out = {1{$random}};
  assign io_VwirePorts_0_18_10_out = {1{$random}};
  assign io_VwirePorts_0_18_11_out = {1{$random}};
  assign io_VwirePorts_0_18_12_out = {1{$random}};
  assign io_VwirePorts_0_18_13_out = {1{$random}};
  assign io_VwirePorts_0_18_14_out = {1{$random}};
  assign io_VwirePorts_0_18_15_out = {1{$random}};
  assign io_VwirePorts_0_19_2_out = {1{$random}};
  assign io_VwirePorts_0_19_6_out = {1{$random}};
  assign io_VwirePorts_0_19_7_out = {1{$random}};
  assign io_VwirePorts_0_19_8_out = {1{$random}};
  assign io_VwirePorts_0_19_9_out = {1{$random}};
  assign io_VwirePorts_0_19_10_out = {1{$random}};
  assign io_VwirePorts_0_19_11_out = {1{$random}};
  assign io_VwirePorts_0_19_12_out = {1{$random}};
  assign io_VwirePorts_0_19_13_out = {1{$random}};
  assign io_VwirePorts_0_19_14_out = {1{$random}};
  assign io_VwirePorts_0_19_15_out = {1{$random}};
  assign io_VwirePorts_0_20_2_out = {1{$random}};
  assign io_VwirePorts_0_20_6_out = {1{$random}};
  assign io_VwirePorts_0_20_7_out = {1{$random}};
  assign io_VwirePorts_0_20_8_out = {1{$random}};
  assign io_VwirePorts_0_20_9_out = {1{$random}};
  assign io_VwirePorts_0_20_10_out = {1{$random}};
  assign io_VwirePorts_0_20_11_out = {1{$random}};
  assign io_VwirePorts_0_20_12_out = {1{$random}};
  assign io_VwirePorts_0_20_13_out = {1{$random}};
  assign io_VwirePorts_0_20_14_out = {1{$random}};
  assign io_VwirePorts_0_20_15_out = {1{$random}};
  assign io_VwirePorts_0_21_2_out = {1{$random}};
  assign io_VwirePorts_0_21_6_out = {1{$random}};
  assign io_VwirePorts_0_21_7_out = {1{$random}};
  assign io_VwirePorts_0_21_8_out = {1{$random}};
  assign io_VwirePorts_0_21_9_out = {1{$random}};
  assign io_VwirePorts_0_21_10_out = {1{$random}};
  assign io_VwirePorts_0_21_11_out = {1{$random}};
  assign io_VwirePorts_0_21_12_out = {1{$random}};
  assign io_VwirePorts_0_21_13_out = {1{$random}};
  assign io_VwirePorts_0_21_14_out = {1{$random}};
  assign io_VwirePorts_0_21_15_out = {1{$random}};
  assign io_VwirePorts_0_22_2_out = {1{$random}};
  assign io_VwirePorts_0_22_6_out = {1{$random}};
  assign io_VwirePorts_0_22_7_out = {1{$random}};
  assign io_VwirePorts_0_22_8_out = {1{$random}};
  assign io_VwirePorts_0_22_9_out = {1{$random}};
  assign io_VwirePorts_0_22_10_out = {1{$random}};
  assign io_VwirePorts_0_22_11_out = {1{$random}};
  assign io_VwirePorts_0_22_12_out = {1{$random}};
  assign io_VwirePorts_0_22_13_out = {1{$random}};
  assign io_VwirePorts_0_22_14_out = {1{$random}};
  assign io_VwirePorts_0_22_15_out = {1{$random}};
  assign io_VwirePorts_1_0_6_out = {1{$random}};
  assign io_VwirePorts_1_0_7_out = {1{$random}};
  assign io_VwirePorts_1_0_8_out = {1{$random}};
  assign io_VwirePorts_1_0_9_out = {1{$random}};
  assign io_VwirePorts_1_0_10_out = {1{$random}};
  assign io_VwirePorts_1_0_11_out = {1{$random}};
  assign io_VwirePorts_1_0_12_out = {1{$random}};
  assign io_VwirePorts_1_0_13_out = {1{$random}};
  assign io_VwirePorts_1_0_14_out = {1{$random}};
  assign io_VwirePorts_1_0_15_out = {1{$random}};
  assign io_VwirePorts_1_1_6_out = {1{$random}};
  assign io_VwirePorts_1_1_7_out = {1{$random}};
  assign io_VwirePorts_1_1_8_out = {1{$random}};
  assign io_VwirePorts_1_1_9_out = {1{$random}};
  assign io_VwirePorts_1_1_10_out = {1{$random}};
  assign io_VwirePorts_1_1_11_out = {1{$random}};
  assign io_VwirePorts_1_1_12_out = {1{$random}};
  assign io_VwirePorts_1_1_13_out = {1{$random}};
  assign io_VwirePorts_1_1_14_out = {1{$random}};
  assign io_VwirePorts_1_1_15_out = {1{$random}};
  assign io_VwirePorts_1_2_6_out = {1{$random}};
  assign io_VwirePorts_1_2_7_out = {1{$random}};
  assign io_VwirePorts_1_2_8_out = {1{$random}};
  assign io_VwirePorts_1_2_9_out = {1{$random}};
  assign io_VwirePorts_1_2_10_out = {1{$random}};
  assign io_VwirePorts_1_2_11_out = {1{$random}};
  assign io_VwirePorts_1_2_12_out = {1{$random}};
  assign io_VwirePorts_1_2_13_out = {1{$random}};
  assign io_VwirePorts_1_2_14_out = {1{$random}};
  assign io_VwirePorts_1_2_15_out = {1{$random}};
  assign io_VwirePorts_1_3_6_out = {1{$random}};
  assign io_VwirePorts_1_3_7_out = {1{$random}};
  assign io_VwirePorts_1_3_8_out = {1{$random}};
  assign io_VwirePorts_1_3_9_out = {1{$random}};
  assign io_VwirePorts_1_3_10_out = {1{$random}};
  assign io_VwirePorts_1_3_11_out = {1{$random}};
  assign io_VwirePorts_1_3_12_out = {1{$random}};
  assign io_VwirePorts_1_3_13_out = {1{$random}};
  assign io_VwirePorts_1_3_14_out = {1{$random}};
  assign io_VwirePorts_1_3_15_out = {1{$random}};
  assign io_VwirePorts_1_4_6_out = {1{$random}};
  assign io_VwirePorts_1_4_7_out = {1{$random}};
  assign io_VwirePorts_1_4_8_out = {1{$random}};
  assign io_VwirePorts_1_4_9_out = {1{$random}};
  assign io_VwirePorts_1_4_10_out = {1{$random}};
  assign io_VwirePorts_1_4_11_out = {1{$random}};
  assign io_VwirePorts_1_4_12_out = {1{$random}};
  assign io_VwirePorts_1_4_13_out = {1{$random}};
  assign io_VwirePorts_1_4_14_out = {1{$random}};
  assign io_VwirePorts_1_4_15_out = {1{$random}};
  assign io_VwirePorts_1_5_6_out = {1{$random}};
  assign io_VwirePorts_1_5_7_out = {1{$random}};
  assign io_VwirePorts_1_5_8_out = {1{$random}};
  assign io_VwirePorts_1_5_9_out = {1{$random}};
  assign io_VwirePorts_1_5_10_out = {1{$random}};
  assign io_VwirePorts_1_5_11_out = {1{$random}};
  assign io_VwirePorts_1_5_12_out = {1{$random}};
  assign io_VwirePorts_1_5_13_out = {1{$random}};
  assign io_VwirePorts_1_5_14_out = {1{$random}};
  assign io_VwirePorts_1_5_15_out = {1{$random}};
  assign io_VwirePorts_1_6_6_out = {1{$random}};
  assign io_VwirePorts_1_6_7_out = {1{$random}};
  assign io_VwirePorts_1_6_8_out = {1{$random}};
  assign io_VwirePorts_1_6_9_out = {1{$random}};
  assign io_VwirePorts_1_6_10_out = {1{$random}};
  assign io_VwirePorts_1_6_11_out = {1{$random}};
  assign io_VwirePorts_1_6_12_out = {1{$random}};
  assign io_VwirePorts_1_6_13_out = {1{$random}};
  assign io_VwirePorts_1_6_14_out = {1{$random}};
  assign io_VwirePorts_1_6_15_out = {1{$random}};
  assign io_VwirePorts_1_7_6_out = {1{$random}};
  assign io_VwirePorts_1_7_7_out = {1{$random}};
  assign io_VwirePorts_1_7_8_out = {1{$random}};
  assign io_VwirePorts_1_7_9_out = {1{$random}};
  assign io_VwirePorts_1_7_10_out = {1{$random}};
  assign io_VwirePorts_1_7_11_out = {1{$random}};
  assign io_VwirePorts_1_7_12_out = {1{$random}};
  assign io_VwirePorts_1_7_13_out = {1{$random}};
  assign io_VwirePorts_1_7_14_out = {1{$random}};
  assign io_VwirePorts_1_7_15_out = {1{$random}};
  assign io_VwirePorts_1_8_6_out = {1{$random}};
  assign io_VwirePorts_1_8_7_out = {1{$random}};
  assign io_VwirePorts_1_8_8_out = {1{$random}};
  assign io_VwirePorts_1_8_9_out = {1{$random}};
  assign io_VwirePorts_1_8_10_out = {1{$random}};
  assign io_VwirePorts_1_8_11_out = {1{$random}};
  assign io_VwirePorts_1_8_12_out = {1{$random}};
  assign io_VwirePorts_1_8_13_out = {1{$random}};
  assign io_VwirePorts_1_8_14_out = {1{$random}};
  assign io_VwirePorts_1_8_15_out = {1{$random}};
  assign io_VwirePorts_1_9_6_out = {1{$random}};
  assign io_VwirePorts_1_9_7_out = {1{$random}};
  assign io_VwirePorts_1_9_8_out = {1{$random}};
  assign io_VwirePorts_1_9_9_out = {1{$random}};
  assign io_VwirePorts_1_9_10_out = {1{$random}};
  assign io_VwirePorts_1_9_11_out = {1{$random}};
  assign io_VwirePorts_1_9_12_out = {1{$random}};
  assign io_VwirePorts_1_9_13_out = {1{$random}};
  assign io_VwirePorts_1_9_14_out = {1{$random}};
  assign io_VwirePorts_1_9_15_out = {1{$random}};
  assign io_VwirePorts_1_10_6_out = {1{$random}};
  assign io_VwirePorts_1_10_7_out = {1{$random}};
  assign io_VwirePorts_1_10_8_out = {1{$random}};
  assign io_VwirePorts_1_10_9_out = {1{$random}};
  assign io_VwirePorts_1_10_10_out = {1{$random}};
  assign io_VwirePorts_1_10_11_out = {1{$random}};
  assign io_VwirePorts_1_10_12_out = {1{$random}};
  assign io_VwirePorts_1_10_13_out = {1{$random}};
  assign io_VwirePorts_1_10_14_out = {1{$random}};
  assign io_VwirePorts_1_10_15_out = {1{$random}};
  assign io_VwirePorts_1_11_6_out = {1{$random}};
  assign io_VwirePorts_1_11_7_out = {1{$random}};
  assign io_VwirePorts_1_11_8_out = {1{$random}};
  assign io_VwirePorts_1_11_9_out = {1{$random}};
  assign io_VwirePorts_1_11_10_out = {1{$random}};
  assign io_VwirePorts_1_11_11_out = {1{$random}};
  assign io_VwirePorts_1_11_12_out = {1{$random}};
  assign io_VwirePorts_1_11_13_out = {1{$random}};
  assign io_VwirePorts_1_11_14_out = {1{$random}};
  assign io_VwirePorts_1_11_15_out = {1{$random}};
  assign io_VwirePorts_1_12_6_out = {1{$random}};
  assign io_VwirePorts_1_12_7_out = {1{$random}};
  assign io_VwirePorts_1_12_8_out = {1{$random}};
  assign io_VwirePorts_1_12_9_out = {1{$random}};
  assign io_VwirePorts_1_12_10_out = {1{$random}};
  assign io_VwirePorts_1_12_11_out = {1{$random}};
  assign io_VwirePorts_1_12_12_out = {1{$random}};
  assign io_VwirePorts_1_12_13_out = {1{$random}};
  assign io_VwirePorts_1_12_14_out = {1{$random}};
  assign io_VwirePorts_1_12_15_out = {1{$random}};
  assign io_VwirePorts_1_13_6_out = {1{$random}};
  assign io_VwirePorts_1_13_7_out = {1{$random}};
  assign io_VwirePorts_1_13_8_out = {1{$random}};
  assign io_VwirePorts_1_13_9_out = {1{$random}};
  assign io_VwirePorts_1_13_10_out = {1{$random}};
  assign io_VwirePorts_1_13_11_out = {1{$random}};
  assign io_VwirePorts_1_13_12_out = {1{$random}};
  assign io_VwirePorts_1_13_13_out = {1{$random}};
  assign io_VwirePorts_1_13_14_out = {1{$random}};
  assign io_VwirePorts_1_13_15_out = {1{$random}};
  assign io_VwirePorts_1_14_6_out = {1{$random}};
  assign io_VwirePorts_1_14_7_out = {1{$random}};
  assign io_VwirePorts_1_14_8_out = {1{$random}};
  assign io_VwirePorts_1_14_9_out = {1{$random}};
  assign io_VwirePorts_1_14_10_out = {1{$random}};
  assign io_VwirePorts_1_14_11_out = {1{$random}};
  assign io_VwirePorts_1_14_12_out = {1{$random}};
  assign io_VwirePorts_1_14_13_out = {1{$random}};
  assign io_VwirePorts_1_14_14_out = {1{$random}};
  assign io_VwirePorts_1_14_15_out = {1{$random}};
  assign io_VwirePorts_1_15_6_out = {1{$random}};
  assign io_VwirePorts_1_15_7_out = {1{$random}};
  assign io_VwirePorts_1_15_8_out = {1{$random}};
  assign io_VwirePorts_1_15_9_out = {1{$random}};
  assign io_VwirePorts_1_15_10_out = {1{$random}};
  assign io_VwirePorts_1_15_11_out = {1{$random}};
  assign io_VwirePorts_1_15_12_out = {1{$random}};
  assign io_VwirePorts_1_15_13_out = {1{$random}};
  assign io_VwirePorts_1_15_14_out = {1{$random}};
  assign io_VwirePorts_1_15_15_out = {1{$random}};
  assign io_VwirePorts_1_16_6_out = {1{$random}};
  assign io_VwirePorts_1_16_7_out = {1{$random}};
  assign io_VwirePorts_1_16_8_out = {1{$random}};
  assign io_VwirePorts_1_16_9_out = {1{$random}};
  assign io_VwirePorts_1_16_10_out = {1{$random}};
  assign io_VwirePorts_1_16_11_out = {1{$random}};
  assign io_VwirePorts_1_16_12_out = {1{$random}};
  assign io_VwirePorts_1_16_13_out = {1{$random}};
  assign io_VwirePorts_1_16_14_out = {1{$random}};
  assign io_VwirePorts_1_16_15_out = {1{$random}};
  assign io_VwirePorts_1_17_6_out = {1{$random}};
  assign io_VwirePorts_1_17_7_out = {1{$random}};
  assign io_VwirePorts_1_17_8_out = {1{$random}};
  assign io_VwirePorts_1_17_9_out = {1{$random}};
  assign io_VwirePorts_1_17_10_out = {1{$random}};
  assign io_VwirePorts_1_17_11_out = {1{$random}};
  assign io_VwirePorts_1_17_12_out = {1{$random}};
  assign io_VwirePorts_1_17_13_out = {1{$random}};
  assign io_VwirePorts_1_17_14_out = {1{$random}};
  assign io_VwirePorts_1_17_15_out = {1{$random}};
  assign io_VwirePorts_1_18_6_out = {1{$random}};
  assign io_VwirePorts_1_18_7_out = {1{$random}};
  assign io_VwirePorts_1_18_8_out = {1{$random}};
  assign io_VwirePorts_1_18_9_out = {1{$random}};
  assign io_VwirePorts_1_18_10_out = {1{$random}};
  assign io_VwirePorts_1_18_11_out = {1{$random}};
  assign io_VwirePorts_1_18_12_out = {1{$random}};
  assign io_VwirePorts_1_18_13_out = {1{$random}};
  assign io_VwirePorts_1_18_14_out = {1{$random}};
  assign io_VwirePorts_1_18_15_out = {1{$random}};
  assign io_VwirePorts_1_19_6_out = {1{$random}};
  assign io_VwirePorts_1_19_7_out = {1{$random}};
  assign io_VwirePorts_1_19_8_out = {1{$random}};
  assign io_VwirePorts_1_19_9_out = {1{$random}};
  assign io_VwirePorts_1_19_10_out = {1{$random}};
  assign io_VwirePorts_1_19_11_out = {1{$random}};
  assign io_VwirePorts_1_19_12_out = {1{$random}};
  assign io_VwirePorts_1_19_13_out = {1{$random}};
  assign io_VwirePorts_1_19_14_out = {1{$random}};
  assign io_VwirePorts_1_19_15_out = {1{$random}};
  assign io_VwirePorts_1_20_6_out = {1{$random}};
  assign io_VwirePorts_1_20_7_out = {1{$random}};
  assign io_VwirePorts_1_20_8_out = {1{$random}};
  assign io_VwirePorts_1_20_9_out = {1{$random}};
  assign io_VwirePorts_1_20_10_out = {1{$random}};
  assign io_VwirePorts_1_20_11_out = {1{$random}};
  assign io_VwirePorts_1_20_12_out = {1{$random}};
  assign io_VwirePorts_1_20_13_out = {1{$random}};
  assign io_VwirePorts_1_20_14_out = {1{$random}};
  assign io_VwirePorts_1_20_15_out = {1{$random}};
  assign io_VwirePorts_1_21_6_out = {1{$random}};
  assign io_VwirePorts_1_21_7_out = {1{$random}};
  assign io_VwirePorts_1_21_8_out = {1{$random}};
  assign io_VwirePorts_1_21_9_out = {1{$random}};
  assign io_VwirePorts_1_21_10_out = {1{$random}};
  assign io_VwirePorts_1_21_11_out = {1{$random}};
  assign io_VwirePorts_1_21_12_out = {1{$random}};
  assign io_VwirePorts_1_21_13_out = {1{$random}};
  assign io_VwirePorts_1_21_14_out = {1{$random}};
  assign io_VwirePorts_1_21_15_out = {1{$random}};
  assign io_VwirePorts_1_22_6_out = {1{$random}};
  assign io_VwirePorts_1_22_7_out = {1{$random}};
  assign io_VwirePorts_1_22_8_out = {1{$random}};
  assign io_VwirePorts_1_22_9_out = {1{$random}};
  assign io_VwirePorts_1_22_10_out = {1{$random}};
  assign io_VwirePorts_1_22_11_out = {1{$random}};
  assign io_VwirePorts_1_22_12_out = {1{$random}};
  assign io_VwirePorts_1_22_13_out = {1{$random}};
  assign io_VwirePorts_1_22_14_out = {1{$random}};
  assign io_VwirePorts_1_22_15_out = {1{$random}};
  assign io_VwirePorts_2_0_6_out = {1{$random}};
  assign io_VwirePorts_2_0_7_out = {1{$random}};
  assign io_VwirePorts_2_0_8_out = {1{$random}};
  assign io_VwirePorts_2_0_9_out = {1{$random}};
  assign io_VwirePorts_2_0_10_out = {1{$random}};
  assign io_VwirePorts_2_0_11_out = {1{$random}};
  assign io_VwirePorts_2_0_12_out = {1{$random}};
  assign io_VwirePorts_2_0_13_out = {1{$random}};
  assign io_VwirePorts_2_0_14_out = {1{$random}};
  assign io_VwirePorts_2_0_15_out = {1{$random}};
  assign io_VwirePorts_2_1_6_out = {1{$random}};
  assign io_VwirePorts_2_1_7_out = {1{$random}};
  assign io_VwirePorts_2_1_8_out = {1{$random}};
  assign io_VwirePorts_2_1_9_out = {1{$random}};
  assign io_VwirePorts_2_1_10_out = {1{$random}};
  assign io_VwirePorts_2_1_11_out = {1{$random}};
  assign io_VwirePorts_2_1_12_out = {1{$random}};
  assign io_VwirePorts_2_1_13_out = {1{$random}};
  assign io_VwirePorts_2_1_14_out = {1{$random}};
  assign io_VwirePorts_2_1_15_out = {1{$random}};
  assign io_VwirePorts_2_2_6_out = {1{$random}};
  assign io_VwirePorts_2_2_7_out = {1{$random}};
  assign io_VwirePorts_2_2_8_out = {1{$random}};
  assign io_VwirePorts_2_2_9_out = {1{$random}};
  assign io_VwirePorts_2_2_10_out = {1{$random}};
  assign io_VwirePorts_2_2_11_out = {1{$random}};
  assign io_VwirePorts_2_2_12_out = {1{$random}};
  assign io_VwirePorts_2_2_13_out = {1{$random}};
  assign io_VwirePorts_2_2_14_out = {1{$random}};
  assign io_VwirePorts_2_2_15_out = {1{$random}};
  assign io_VwirePorts_2_3_6_out = {1{$random}};
  assign io_VwirePorts_2_3_7_out = {1{$random}};
  assign io_VwirePorts_2_3_8_out = {1{$random}};
  assign io_VwirePorts_2_3_9_out = {1{$random}};
  assign io_VwirePorts_2_3_10_out = {1{$random}};
  assign io_VwirePorts_2_3_11_out = {1{$random}};
  assign io_VwirePorts_2_3_12_out = {1{$random}};
  assign io_VwirePorts_2_3_13_out = {1{$random}};
  assign io_VwirePorts_2_3_14_out = {1{$random}};
  assign io_VwirePorts_2_3_15_out = {1{$random}};
  assign io_VwirePorts_2_4_6_out = {1{$random}};
  assign io_VwirePorts_2_4_7_out = {1{$random}};
  assign io_VwirePorts_2_4_8_out = {1{$random}};
  assign io_VwirePorts_2_4_9_out = {1{$random}};
  assign io_VwirePorts_2_4_10_out = {1{$random}};
  assign io_VwirePorts_2_4_11_out = {1{$random}};
  assign io_VwirePorts_2_4_12_out = {1{$random}};
  assign io_VwirePorts_2_4_13_out = {1{$random}};
  assign io_VwirePorts_2_4_14_out = {1{$random}};
  assign io_VwirePorts_2_4_15_out = {1{$random}};
  assign io_VwirePorts_2_5_6_out = {1{$random}};
  assign io_VwirePorts_2_5_7_out = {1{$random}};
  assign io_VwirePorts_2_5_8_out = {1{$random}};
  assign io_VwirePorts_2_5_9_out = {1{$random}};
  assign io_VwirePorts_2_5_10_out = {1{$random}};
  assign io_VwirePorts_2_5_11_out = {1{$random}};
  assign io_VwirePorts_2_5_12_out = {1{$random}};
  assign io_VwirePorts_2_5_13_out = {1{$random}};
  assign io_VwirePorts_2_5_14_out = {1{$random}};
  assign io_VwirePorts_2_5_15_out = {1{$random}};
  assign io_VwirePorts_2_6_6_out = {1{$random}};
  assign io_VwirePorts_2_6_7_out = {1{$random}};
  assign io_VwirePorts_2_6_8_out = {1{$random}};
  assign io_VwirePorts_2_6_9_out = {1{$random}};
  assign io_VwirePorts_2_6_10_out = {1{$random}};
  assign io_VwirePorts_2_6_11_out = {1{$random}};
  assign io_VwirePorts_2_6_12_out = {1{$random}};
  assign io_VwirePorts_2_6_13_out = {1{$random}};
  assign io_VwirePorts_2_6_14_out = {1{$random}};
  assign io_VwirePorts_2_6_15_out = {1{$random}};
  assign io_VwirePorts_2_7_6_out = {1{$random}};
  assign io_VwirePorts_2_7_7_out = {1{$random}};
  assign io_VwirePorts_2_7_8_out = {1{$random}};
  assign io_VwirePorts_2_7_9_out = {1{$random}};
  assign io_VwirePorts_2_7_10_out = {1{$random}};
  assign io_VwirePorts_2_7_11_out = {1{$random}};
  assign io_VwirePorts_2_7_12_out = {1{$random}};
  assign io_VwirePorts_2_7_13_out = {1{$random}};
  assign io_VwirePorts_2_7_14_out = {1{$random}};
  assign io_VwirePorts_2_7_15_out = {1{$random}};
  assign io_VwirePorts_2_8_6_out = {1{$random}};
  assign io_VwirePorts_2_8_7_out = {1{$random}};
  assign io_VwirePorts_2_8_8_out = {1{$random}};
  assign io_VwirePorts_2_8_9_out = {1{$random}};
  assign io_VwirePorts_2_8_10_out = {1{$random}};
  assign io_VwirePorts_2_8_11_out = {1{$random}};
  assign io_VwirePorts_2_8_12_out = {1{$random}};
  assign io_VwirePorts_2_8_13_out = {1{$random}};
  assign io_VwirePorts_2_8_14_out = {1{$random}};
  assign io_VwirePorts_2_8_15_out = {1{$random}};
  assign io_VwirePorts_2_9_6_out = {1{$random}};
  assign io_VwirePorts_2_9_7_out = {1{$random}};
  assign io_VwirePorts_2_9_8_out = {1{$random}};
  assign io_VwirePorts_2_9_9_out = {1{$random}};
  assign io_VwirePorts_2_9_10_out = {1{$random}};
  assign io_VwirePorts_2_9_11_out = {1{$random}};
  assign io_VwirePorts_2_9_12_out = {1{$random}};
  assign io_VwirePorts_2_9_13_out = {1{$random}};
  assign io_VwirePorts_2_9_14_out = {1{$random}};
  assign io_VwirePorts_2_9_15_out = {1{$random}};
  assign io_VwirePorts_2_10_6_out = {1{$random}};
  assign io_VwirePorts_2_10_7_out = {1{$random}};
  assign io_VwirePorts_2_10_8_out = {1{$random}};
  assign io_VwirePorts_2_10_9_out = {1{$random}};
  assign io_VwirePorts_2_10_10_out = {1{$random}};
  assign io_VwirePorts_2_10_11_out = {1{$random}};
  assign io_VwirePorts_2_10_12_out = {1{$random}};
  assign io_VwirePorts_2_10_13_out = {1{$random}};
  assign io_VwirePorts_2_10_14_out = {1{$random}};
  assign io_VwirePorts_2_10_15_out = {1{$random}};
  assign io_VwirePorts_2_11_6_out = {1{$random}};
  assign io_VwirePorts_2_11_7_out = {1{$random}};
  assign io_VwirePorts_2_11_8_out = {1{$random}};
  assign io_VwirePorts_2_11_9_out = {1{$random}};
  assign io_VwirePorts_2_11_10_out = {1{$random}};
  assign io_VwirePorts_2_11_11_out = {1{$random}};
  assign io_VwirePorts_2_11_12_out = {1{$random}};
  assign io_VwirePorts_2_11_13_out = {1{$random}};
  assign io_VwirePorts_2_11_14_out = {1{$random}};
  assign io_VwirePorts_2_11_15_out = {1{$random}};
  assign io_VwirePorts_2_12_6_out = {1{$random}};
  assign io_VwirePorts_2_12_7_out = {1{$random}};
  assign io_VwirePorts_2_12_8_out = {1{$random}};
  assign io_VwirePorts_2_12_9_out = {1{$random}};
  assign io_VwirePorts_2_12_10_out = {1{$random}};
  assign io_VwirePorts_2_12_11_out = {1{$random}};
  assign io_VwirePorts_2_12_12_out = {1{$random}};
  assign io_VwirePorts_2_12_13_out = {1{$random}};
  assign io_VwirePorts_2_12_14_out = {1{$random}};
  assign io_VwirePorts_2_12_15_out = {1{$random}};
  assign io_VwirePorts_2_13_6_out = {1{$random}};
  assign io_VwirePorts_2_13_7_out = {1{$random}};
  assign io_VwirePorts_2_13_8_out = {1{$random}};
  assign io_VwirePorts_2_13_9_out = {1{$random}};
  assign io_VwirePorts_2_13_10_out = {1{$random}};
  assign io_VwirePorts_2_13_11_out = {1{$random}};
  assign io_VwirePorts_2_13_12_out = {1{$random}};
  assign io_VwirePorts_2_13_13_out = {1{$random}};
  assign io_VwirePorts_2_13_14_out = {1{$random}};
  assign io_VwirePorts_2_13_15_out = {1{$random}};
  assign io_VwirePorts_2_14_6_out = {1{$random}};
  assign io_VwirePorts_2_14_7_out = {1{$random}};
  assign io_VwirePorts_2_14_8_out = {1{$random}};
  assign io_VwirePorts_2_14_9_out = {1{$random}};
  assign io_VwirePorts_2_14_10_out = {1{$random}};
  assign io_VwirePorts_2_14_11_out = {1{$random}};
  assign io_VwirePorts_2_14_12_out = {1{$random}};
  assign io_VwirePorts_2_14_13_out = {1{$random}};
  assign io_VwirePorts_2_14_14_out = {1{$random}};
  assign io_VwirePorts_2_14_15_out = {1{$random}};
  assign io_VwirePorts_2_15_6_out = {1{$random}};
  assign io_VwirePorts_2_15_7_out = {1{$random}};
  assign io_VwirePorts_2_15_8_out = {1{$random}};
  assign io_VwirePorts_2_15_9_out = {1{$random}};
  assign io_VwirePorts_2_15_10_out = {1{$random}};
  assign io_VwirePorts_2_15_11_out = {1{$random}};
  assign io_VwirePorts_2_15_12_out = {1{$random}};
  assign io_VwirePorts_2_15_13_out = {1{$random}};
  assign io_VwirePorts_2_15_14_out = {1{$random}};
  assign io_VwirePorts_2_15_15_out = {1{$random}};
  assign io_VwirePorts_2_16_6_out = {1{$random}};
  assign io_VwirePorts_2_16_7_out = {1{$random}};
  assign io_VwirePorts_2_16_8_out = {1{$random}};
  assign io_VwirePorts_2_16_9_out = {1{$random}};
  assign io_VwirePorts_2_16_10_out = {1{$random}};
  assign io_VwirePorts_2_16_11_out = {1{$random}};
  assign io_VwirePorts_2_16_12_out = {1{$random}};
  assign io_VwirePorts_2_16_13_out = {1{$random}};
  assign io_VwirePorts_2_16_14_out = {1{$random}};
  assign io_VwirePorts_2_16_15_out = {1{$random}};
  assign io_VwirePorts_2_17_6_out = {1{$random}};
  assign io_VwirePorts_2_17_7_out = {1{$random}};
  assign io_VwirePorts_2_17_8_out = {1{$random}};
  assign io_VwirePorts_2_17_9_out = {1{$random}};
  assign io_VwirePorts_2_17_10_out = {1{$random}};
  assign io_VwirePorts_2_17_11_out = {1{$random}};
  assign io_VwirePorts_2_17_12_out = {1{$random}};
  assign io_VwirePorts_2_17_13_out = {1{$random}};
  assign io_VwirePorts_2_17_14_out = {1{$random}};
  assign io_VwirePorts_2_17_15_out = {1{$random}};
  assign io_VwirePorts_2_18_6_out = {1{$random}};
  assign io_VwirePorts_2_18_7_out = {1{$random}};
  assign io_VwirePorts_2_18_8_out = {1{$random}};
  assign io_VwirePorts_2_18_9_out = {1{$random}};
  assign io_VwirePorts_2_18_10_out = {1{$random}};
  assign io_VwirePorts_2_18_11_out = {1{$random}};
  assign io_VwirePorts_2_18_12_out = {1{$random}};
  assign io_VwirePorts_2_18_13_out = {1{$random}};
  assign io_VwirePorts_2_18_14_out = {1{$random}};
  assign io_VwirePorts_2_18_15_out = {1{$random}};
  assign io_VwirePorts_2_19_6_out = {1{$random}};
  assign io_VwirePorts_2_19_7_out = {1{$random}};
  assign io_VwirePorts_2_19_8_out = {1{$random}};
  assign io_VwirePorts_2_19_9_out = {1{$random}};
  assign io_VwirePorts_2_19_10_out = {1{$random}};
  assign io_VwirePorts_2_19_11_out = {1{$random}};
  assign io_VwirePorts_2_19_12_out = {1{$random}};
  assign io_VwirePorts_2_19_13_out = {1{$random}};
  assign io_VwirePorts_2_19_14_out = {1{$random}};
  assign io_VwirePorts_2_19_15_out = {1{$random}};
  assign io_VwirePorts_2_20_6_out = {1{$random}};
  assign io_VwirePorts_2_20_7_out = {1{$random}};
  assign io_VwirePorts_2_20_8_out = {1{$random}};
  assign io_VwirePorts_2_20_9_out = {1{$random}};
  assign io_VwirePorts_2_20_10_out = {1{$random}};
  assign io_VwirePorts_2_20_11_out = {1{$random}};
  assign io_VwirePorts_2_20_12_out = {1{$random}};
  assign io_VwirePorts_2_20_13_out = {1{$random}};
  assign io_VwirePorts_2_20_14_out = {1{$random}};
  assign io_VwirePorts_2_20_15_out = {1{$random}};
  assign io_VwirePorts_2_21_6_out = {1{$random}};
  assign io_VwirePorts_2_21_7_out = {1{$random}};
  assign io_VwirePorts_2_21_8_out = {1{$random}};
  assign io_VwirePorts_2_21_9_out = {1{$random}};
  assign io_VwirePorts_2_21_10_out = {1{$random}};
  assign io_VwirePorts_2_21_11_out = {1{$random}};
  assign io_VwirePorts_2_21_12_out = {1{$random}};
  assign io_VwirePorts_2_21_13_out = {1{$random}};
  assign io_VwirePorts_2_21_14_out = {1{$random}};
  assign io_VwirePorts_2_21_15_out = {1{$random}};
  assign io_VwirePorts_2_22_6_out = {1{$random}};
  assign io_VwirePorts_2_22_7_out = {1{$random}};
  assign io_VwirePorts_2_22_8_out = {1{$random}};
  assign io_VwirePorts_2_22_9_out = {1{$random}};
  assign io_VwirePorts_2_22_10_out = {1{$random}};
  assign io_VwirePorts_2_22_11_out = {1{$random}};
  assign io_VwirePorts_2_22_12_out = {1{$random}};
  assign io_VwirePorts_2_22_13_out = {1{$random}};
  assign io_VwirePorts_2_22_14_out = {1{$random}};
  assign io_VwirePorts_2_22_15_out = {1{$random}};
  assign io_VwirePorts_3_0_2_out = {1{$random}};
  assign io_VwirePorts_3_0_6_out = {1{$random}};
  assign io_VwirePorts_3_0_7_out = {1{$random}};
  assign io_VwirePorts_3_0_8_out = {1{$random}};
  assign io_VwirePorts_3_0_9_out = {1{$random}};
  assign io_VwirePorts_3_0_10_out = {1{$random}};
  assign io_VwirePorts_3_0_11_out = {1{$random}};
  assign io_VwirePorts_3_0_12_out = {1{$random}};
  assign io_VwirePorts_3_0_13_out = {1{$random}};
  assign io_VwirePorts_3_0_14_out = {1{$random}};
  assign io_VwirePorts_3_0_15_out = {1{$random}};
  assign io_VwirePorts_3_1_2_out = {1{$random}};
  assign io_VwirePorts_3_1_6_out = {1{$random}};
  assign io_VwirePorts_3_1_7_out = {1{$random}};
  assign io_VwirePorts_3_1_8_out = {1{$random}};
  assign io_VwirePorts_3_1_9_out = {1{$random}};
  assign io_VwirePorts_3_1_10_out = {1{$random}};
  assign io_VwirePorts_3_1_11_out = {1{$random}};
  assign io_VwirePorts_3_1_12_out = {1{$random}};
  assign io_VwirePorts_3_1_13_out = {1{$random}};
  assign io_VwirePorts_3_1_14_out = {1{$random}};
  assign io_VwirePorts_3_1_15_out = {1{$random}};
  assign io_VwirePorts_3_2_2_out = {1{$random}};
  assign io_VwirePorts_3_2_6_out = {1{$random}};
  assign io_VwirePorts_3_2_7_out = {1{$random}};
  assign io_VwirePorts_3_2_8_out = {1{$random}};
  assign io_VwirePorts_3_2_9_out = {1{$random}};
  assign io_VwirePorts_3_2_10_out = {1{$random}};
  assign io_VwirePorts_3_2_11_out = {1{$random}};
  assign io_VwirePorts_3_2_12_out = {1{$random}};
  assign io_VwirePorts_3_2_13_out = {1{$random}};
  assign io_VwirePorts_3_2_14_out = {1{$random}};
  assign io_VwirePorts_3_2_15_out = {1{$random}};
  assign io_VwirePorts_3_3_2_out = {1{$random}};
  assign io_VwirePorts_3_3_6_out = {1{$random}};
  assign io_VwirePorts_3_3_7_out = {1{$random}};
  assign io_VwirePorts_3_3_8_out = {1{$random}};
  assign io_VwirePorts_3_3_9_out = {1{$random}};
  assign io_VwirePorts_3_3_10_out = {1{$random}};
  assign io_VwirePorts_3_3_11_out = {1{$random}};
  assign io_VwirePorts_3_3_12_out = {1{$random}};
  assign io_VwirePorts_3_3_13_out = {1{$random}};
  assign io_VwirePorts_3_3_14_out = {1{$random}};
  assign io_VwirePorts_3_3_15_out = {1{$random}};
  assign io_VwirePorts_3_4_2_out = {1{$random}};
  assign io_VwirePorts_3_4_6_out = {1{$random}};
  assign io_VwirePorts_3_4_7_out = {1{$random}};
  assign io_VwirePorts_3_4_8_out = {1{$random}};
  assign io_VwirePorts_3_4_9_out = {1{$random}};
  assign io_VwirePorts_3_4_10_out = {1{$random}};
  assign io_VwirePorts_3_4_11_out = {1{$random}};
  assign io_VwirePorts_3_4_12_out = {1{$random}};
  assign io_VwirePorts_3_4_13_out = {1{$random}};
  assign io_VwirePorts_3_4_14_out = {1{$random}};
  assign io_VwirePorts_3_4_15_out = {1{$random}};
  assign io_VwirePorts_3_5_2_out = {1{$random}};
  assign io_VwirePorts_3_5_6_out = {1{$random}};
  assign io_VwirePorts_3_5_7_out = {1{$random}};
  assign io_VwirePorts_3_5_8_out = {1{$random}};
  assign io_VwirePorts_3_5_9_out = {1{$random}};
  assign io_VwirePorts_3_5_10_out = {1{$random}};
  assign io_VwirePorts_3_5_11_out = {1{$random}};
  assign io_VwirePorts_3_5_12_out = {1{$random}};
  assign io_VwirePorts_3_5_13_out = {1{$random}};
  assign io_VwirePorts_3_5_14_out = {1{$random}};
  assign io_VwirePorts_3_5_15_out = {1{$random}};
  assign io_VwirePorts_3_6_2_out = {1{$random}};
  assign io_VwirePorts_3_6_6_out = {1{$random}};
  assign io_VwirePorts_3_6_7_out = {1{$random}};
  assign io_VwirePorts_3_6_8_out = {1{$random}};
  assign io_VwirePorts_3_6_9_out = {1{$random}};
  assign io_VwirePorts_3_6_10_out = {1{$random}};
  assign io_VwirePorts_3_6_11_out = {1{$random}};
  assign io_VwirePorts_3_6_12_out = {1{$random}};
  assign io_VwirePorts_3_6_13_out = {1{$random}};
  assign io_VwirePorts_3_6_14_out = {1{$random}};
  assign io_VwirePorts_3_6_15_out = {1{$random}};
  assign io_VwirePorts_3_7_2_out = {1{$random}};
  assign io_VwirePorts_3_7_6_out = {1{$random}};
  assign io_VwirePorts_3_7_7_out = {1{$random}};
  assign io_VwirePorts_3_7_8_out = {1{$random}};
  assign io_VwirePorts_3_7_9_out = {1{$random}};
  assign io_VwirePorts_3_7_10_out = {1{$random}};
  assign io_VwirePorts_3_7_11_out = {1{$random}};
  assign io_VwirePorts_3_7_12_out = {1{$random}};
  assign io_VwirePorts_3_7_13_out = {1{$random}};
  assign io_VwirePorts_3_7_14_out = {1{$random}};
  assign io_VwirePorts_3_7_15_out = {1{$random}};
  assign io_VwirePorts_3_8_2_out = {1{$random}};
  assign io_VwirePorts_3_8_6_out = {1{$random}};
  assign io_VwirePorts_3_8_7_out = {1{$random}};
  assign io_VwirePorts_3_8_8_out = {1{$random}};
  assign io_VwirePorts_3_8_9_out = {1{$random}};
  assign io_VwirePorts_3_8_10_out = {1{$random}};
  assign io_VwirePorts_3_8_11_out = {1{$random}};
  assign io_VwirePorts_3_8_12_out = {1{$random}};
  assign io_VwirePorts_3_8_13_out = {1{$random}};
  assign io_VwirePorts_3_8_14_out = {1{$random}};
  assign io_VwirePorts_3_8_15_out = {1{$random}};
  assign io_VwirePorts_3_9_2_out = {1{$random}};
  assign io_VwirePorts_3_9_6_out = {1{$random}};
  assign io_VwirePorts_3_9_7_out = {1{$random}};
  assign io_VwirePorts_3_9_8_out = {1{$random}};
  assign io_VwirePorts_3_9_9_out = {1{$random}};
  assign io_VwirePorts_3_9_10_out = {1{$random}};
  assign io_VwirePorts_3_9_11_out = {1{$random}};
  assign io_VwirePorts_3_9_12_out = {1{$random}};
  assign io_VwirePorts_3_9_13_out = {1{$random}};
  assign io_VwirePorts_3_9_14_out = {1{$random}};
  assign io_VwirePorts_3_9_15_out = {1{$random}};
  assign io_VwirePorts_3_10_2_out = {1{$random}};
  assign io_VwirePorts_3_10_6_out = {1{$random}};
  assign io_VwirePorts_3_10_7_out = {1{$random}};
  assign io_VwirePorts_3_10_8_out = {1{$random}};
  assign io_VwirePorts_3_10_9_out = {1{$random}};
  assign io_VwirePorts_3_10_10_out = {1{$random}};
  assign io_VwirePorts_3_10_11_out = {1{$random}};
  assign io_VwirePorts_3_10_12_out = {1{$random}};
  assign io_VwirePorts_3_10_13_out = {1{$random}};
  assign io_VwirePorts_3_10_14_out = {1{$random}};
  assign io_VwirePorts_3_10_15_out = {1{$random}};
  assign io_VwirePorts_3_11_2_out = {1{$random}};
  assign io_VwirePorts_3_11_6_out = {1{$random}};
  assign io_VwirePorts_3_11_7_out = {1{$random}};
  assign io_VwirePorts_3_11_8_out = {1{$random}};
  assign io_VwirePorts_3_11_9_out = {1{$random}};
  assign io_VwirePorts_3_11_10_out = {1{$random}};
  assign io_VwirePorts_3_11_11_out = {1{$random}};
  assign io_VwirePorts_3_11_12_out = {1{$random}};
  assign io_VwirePorts_3_11_13_out = {1{$random}};
  assign io_VwirePorts_3_11_14_out = {1{$random}};
  assign io_VwirePorts_3_11_15_out = {1{$random}};
  assign io_VwirePorts_3_12_2_out = {1{$random}};
  assign io_VwirePorts_3_12_6_out = {1{$random}};
  assign io_VwirePorts_3_12_7_out = {1{$random}};
  assign io_VwirePorts_3_12_8_out = {1{$random}};
  assign io_VwirePorts_3_12_9_out = {1{$random}};
  assign io_VwirePorts_3_12_10_out = {1{$random}};
  assign io_VwirePorts_3_12_11_out = {1{$random}};
  assign io_VwirePorts_3_12_12_out = {1{$random}};
  assign io_VwirePorts_3_12_13_out = {1{$random}};
  assign io_VwirePorts_3_12_14_out = {1{$random}};
  assign io_VwirePorts_3_12_15_out = {1{$random}};
  assign io_VwirePorts_3_13_2_out = {1{$random}};
  assign io_VwirePorts_3_13_6_out = {1{$random}};
  assign io_VwirePorts_3_13_7_out = {1{$random}};
  assign io_VwirePorts_3_13_8_out = {1{$random}};
  assign io_VwirePorts_3_13_9_out = {1{$random}};
  assign io_VwirePorts_3_13_10_out = {1{$random}};
  assign io_VwirePorts_3_13_11_out = {1{$random}};
  assign io_VwirePorts_3_13_12_out = {1{$random}};
  assign io_VwirePorts_3_13_13_out = {1{$random}};
  assign io_VwirePorts_3_13_14_out = {1{$random}};
  assign io_VwirePorts_3_13_15_out = {1{$random}};
  assign io_VwirePorts_3_14_2_out = {1{$random}};
  assign io_VwirePorts_3_14_6_out = {1{$random}};
  assign io_VwirePorts_3_14_7_out = {1{$random}};
  assign io_VwirePorts_3_14_8_out = {1{$random}};
  assign io_VwirePorts_3_14_9_out = {1{$random}};
  assign io_VwirePorts_3_14_10_out = {1{$random}};
  assign io_VwirePorts_3_14_11_out = {1{$random}};
  assign io_VwirePorts_3_14_12_out = {1{$random}};
  assign io_VwirePorts_3_14_13_out = {1{$random}};
  assign io_VwirePorts_3_14_14_out = {1{$random}};
  assign io_VwirePorts_3_14_15_out = {1{$random}};
  assign io_VwirePorts_3_15_2_out = {1{$random}};
  assign io_VwirePorts_3_15_6_out = {1{$random}};
  assign io_VwirePorts_3_15_7_out = {1{$random}};
  assign io_VwirePorts_3_15_8_out = {1{$random}};
  assign io_VwirePorts_3_15_9_out = {1{$random}};
  assign io_VwirePorts_3_15_10_out = {1{$random}};
  assign io_VwirePorts_3_15_11_out = {1{$random}};
  assign io_VwirePorts_3_15_12_out = {1{$random}};
  assign io_VwirePorts_3_15_13_out = {1{$random}};
  assign io_VwirePorts_3_15_14_out = {1{$random}};
  assign io_VwirePorts_3_15_15_out = {1{$random}};
  assign io_VwirePorts_3_16_2_out = {1{$random}};
  assign io_VwirePorts_3_16_6_out = {1{$random}};
  assign io_VwirePorts_3_16_7_out = {1{$random}};
  assign io_VwirePorts_3_16_8_out = {1{$random}};
  assign io_VwirePorts_3_16_9_out = {1{$random}};
  assign io_VwirePorts_3_16_10_out = {1{$random}};
  assign io_VwirePorts_3_16_11_out = {1{$random}};
  assign io_VwirePorts_3_16_12_out = {1{$random}};
  assign io_VwirePorts_3_16_13_out = {1{$random}};
  assign io_VwirePorts_3_16_14_out = {1{$random}};
  assign io_VwirePorts_3_16_15_out = {1{$random}};
  assign io_VwirePorts_3_17_2_out = {1{$random}};
  assign io_VwirePorts_3_17_6_out = {1{$random}};
  assign io_VwirePorts_3_17_7_out = {1{$random}};
  assign io_VwirePorts_3_17_8_out = {1{$random}};
  assign io_VwirePorts_3_17_9_out = {1{$random}};
  assign io_VwirePorts_3_17_10_out = {1{$random}};
  assign io_VwirePorts_3_17_11_out = {1{$random}};
  assign io_VwirePorts_3_17_12_out = {1{$random}};
  assign io_VwirePorts_3_17_13_out = {1{$random}};
  assign io_VwirePorts_3_17_14_out = {1{$random}};
  assign io_VwirePorts_3_17_15_out = {1{$random}};
  assign io_VwirePorts_3_18_2_out = {1{$random}};
  assign io_VwirePorts_3_18_6_out = {1{$random}};
  assign io_VwirePorts_3_18_7_out = {1{$random}};
  assign io_VwirePorts_3_18_8_out = {1{$random}};
  assign io_VwirePorts_3_18_9_out = {1{$random}};
  assign io_VwirePorts_3_18_10_out = {1{$random}};
  assign io_VwirePorts_3_18_11_out = {1{$random}};
  assign io_VwirePorts_3_18_12_out = {1{$random}};
  assign io_VwirePorts_3_18_13_out = {1{$random}};
  assign io_VwirePorts_3_18_14_out = {1{$random}};
  assign io_VwirePorts_3_18_15_out = {1{$random}};
  assign io_VwirePorts_3_19_2_out = {1{$random}};
  assign io_VwirePorts_3_19_6_out = {1{$random}};
  assign io_VwirePorts_3_19_7_out = {1{$random}};
  assign io_VwirePorts_3_19_8_out = {1{$random}};
  assign io_VwirePorts_3_19_9_out = {1{$random}};
  assign io_VwirePorts_3_19_10_out = {1{$random}};
  assign io_VwirePorts_3_19_11_out = {1{$random}};
  assign io_VwirePorts_3_19_12_out = {1{$random}};
  assign io_VwirePorts_3_19_13_out = {1{$random}};
  assign io_VwirePorts_3_19_14_out = {1{$random}};
  assign io_VwirePorts_3_19_15_out = {1{$random}};
  assign io_VwirePorts_3_20_2_out = {1{$random}};
  assign io_VwirePorts_3_20_6_out = {1{$random}};
  assign io_VwirePorts_3_20_7_out = {1{$random}};
  assign io_VwirePorts_3_20_8_out = {1{$random}};
  assign io_VwirePorts_3_20_9_out = {1{$random}};
  assign io_VwirePorts_3_20_10_out = {1{$random}};
  assign io_VwirePorts_3_20_11_out = {1{$random}};
  assign io_VwirePorts_3_20_12_out = {1{$random}};
  assign io_VwirePorts_3_20_13_out = {1{$random}};
  assign io_VwirePorts_3_20_14_out = {1{$random}};
  assign io_VwirePorts_3_20_15_out = {1{$random}};
  assign io_VwirePorts_3_21_2_out = {1{$random}};
  assign io_VwirePorts_3_21_6_out = {1{$random}};
  assign io_VwirePorts_3_21_7_out = {1{$random}};
  assign io_VwirePorts_3_21_8_out = {1{$random}};
  assign io_VwirePorts_3_21_9_out = {1{$random}};
  assign io_VwirePorts_3_21_10_out = {1{$random}};
  assign io_VwirePorts_3_21_11_out = {1{$random}};
  assign io_VwirePorts_3_21_12_out = {1{$random}};
  assign io_VwirePorts_3_21_13_out = {1{$random}};
  assign io_VwirePorts_3_21_14_out = {1{$random}};
  assign io_VwirePorts_3_21_15_out = {1{$random}};
  assign io_VwirePorts_3_22_2_out = {1{$random}};
  assign io_VwirePorts_3_22_6_out = {1{$random}};
  assign io_VwirePorts_3_22_7_out = {1{$random}};
  assign io_VwirePorts_3_22_8_out = {1{$random}};
  assign io_VwirePorts_3_22_9_out = {1{$random}};
  assign io_VwirePorts_3_22_10_out = {1{$random}};
  assign io_VwirePorts_3_22_11_out = {1{$random}};
  assign io_VwirePorts_3_22_12_out = {1{$random}};
  assign io_VwirePorts_3_22_13_out = {1{$random}};
  assign io_VwirePorts_3_22_14_out = {1{$random}};
  assign io_VwirePorts_3_22_15_out = {1{$random}};
// synthesis translate_on
`endif
  assign io_VwirePorts_0_0_0_out = Vwire_138_io_out;
  assign io_VwirePorts_0_0_1_out = Vwire_23_io_out;
  assign io_VwirePorts_0_0_3_out = Vwire_115_io_out;
  assign io_VwirePorts_0_0_4_out = Vwire_69_io_out;
  assign io_VwirePorts_0_0_5_out = Vwire_161_io_out;
  assign io_VwirePorts_0_1_0_out = Vwire_139_io_out;
  assign io_VwirePorts_0_1_1_out = Vwire_24_io_out;
  assign io_VwirePorts_0_1_3_out = Vwire_116_io_out;
  assign io_VwirePorts_0_1_4_out = Vwire_70_io_out;
  assign io_VwirePorts_0_1_5_out = Vwire_162_io_out;
  assign io_VwirePorts_0_2_0_out = Vwire_140_io_out;
  assign io_VwirePorts_0_2_1_out = Vwire_25_io_out;
  assign io_VwirePorts_0_2_3_out = Vwire_117_io_out;
  assign io_VwirePorts_0_2_4_out = Vwire_71_io_out;
  assign io_VwirePorts_0_2_5_out = Vwire_163_io_out;
  assign io_VwirePorts_0_3_0_out = Vwire_141_io_out;
  assign io_VwirePorts_0_3_1_out = Vwire_26_io_out;
  assign io_VwirePorts_0_3_3_out = Vwire_118_io_out;
  assign io_VwirePorts_0_3_4_out = Vwire_72_io_out;
  assign io_VwirePorts_0_3_5_out = Vwire_164_io_out;
  assign io_VwirePorts_0_4_0_out = Vwire_142_io_out;
  assign io_VwirePorts_0_4_1_out = Vwire_27_io_out;
  assign io_VwirePorts_0_4_3_out = Vwire_119_io_out;
  assign io_VwirePorts_0_4_4_out = Vwire_73_io_out;
  assign io_VwirePorts_0_4_5_out = Vwire_165_io_out;
  assign io_VwirePorts_0_5_0_out = Vwire_143_io_out;
  assign io_VwirePorts_0_5_1_out = Vwire_28_io_out;
  assign io_VwirePorts_0_5_3_out = Vwire_120_io_out;
  assign io_VwirePorts_0_5_4_out = Vwire_74_io_out;
  assign io_VwirePorts_0_5_5_out = Vwire_166_io_out;
  assign io_VwirePorts_0_6_0_out = Vwire_144_io_out;
  assign io_VwirePorts_0_6_1_out = Vwire_29_io_out;
  assign io_VwirePorts_0_6_3_out = Vwire_121_io_out;
  assign io_VwirePorts_0_6_4_out = Vwire_75_io_out;
  assign io_VwirePorts_0_6_5_out = Vwire_167_io_out;
  assign io_VwirePorts_0_7_0_out = Vwire_145_io_out;
  assign io_VwirePorts_0_7_1_out = Vwire_30_io_out;
  assign io_VwirePorts_0_7_3_out = Vwire_122_io_out;
  assign io_VwirePorts_0_7_4_out = Vwire_76_io_out;
  assign io_VwirePorts_0_7_5_out = Vwire_168_io_out;
  assign io_VwirePorts_0_8_0_out = Vwire_146_io_out;
  assign io_VwirePorts_0_8_1_out = Vwire_31_io_out;
  assign io_VwirePorts_0_8_3_out = Vwire_123_io_out;
  assign io_VwirePorts_0_8_4_out = Vwire_77_io_out;
  assign io_VwirePorts_0_8_5_out = Vwire_169_io_out;
  assign io_VwirePorts_0_9_0_out = Vwire_147_io_out;
  assign io_VwirePorts_0_9_1_out = Vwire_32_io_out;
  assign io_VwirePorts_0_9_3_out = Vwire_124_io_out;
  assign io_VwirePorts_0_9_4_out = Vwire_78_io_out;
  assign io_VwirePorts_0_9_5_out = Vwire_170_io_out;
  assign io_VwirePorts_0_10_0_out = Vwire_148_io_out;
  assign io_VwirePorts_0_10_1_out = Vwire_33_io_out;
  assign io_VwirePorts_0_10_3_out = Vwire_125_io_out;
  assign io_VwirePorts_0_10_4_out = Vwire_79_io_out;
  assign io_VwirePorts_0_10_5_out = Vwire_171_io_out;
  assign io_VwirePorts_0_11_0_out = Vwire_149_io_out;
  assign io_VwirePorts_0_11_1_out = Vwire_34_io_out;
  assign io_VwirePorts_0_11_3_out = Vwire_126_io_out;
  assign io_VwirePorts_0_11_4_out = Vwire_80_io_out;
  assign io_VwirePorts_0_11_5_out = Vwire_172_io_out;
  assign io_VwirePorts_0_12_0_out = Vwire_150_io_out;
  assign io_VwirePorts_0_12_1_out = Vwire_35_io_out;
  assign io_VwirePorts_0_12_3_out = Vwire_127_io_out;
  assign io_VwirePorts_0_12_4_out = Vwire_81_io_out;
  assign io_VwirePorts_0_12_5_out = Vwire_173_io_out;
  assign io_VwirePorts_0_13_0_out = Vwire_151_io_out;
  assign io_VwirePorts_0_13_1_out = Vwire_36_io_out;
  assign io_VwirePorts_0_13_3_out = Vwire_128_io_out;
  assign io_VwirePorts_0_13_4_out = Vwire_82_io_out;
  assign io_VwirePorts_0_13_5_out = Vwire_174_io_out;
  assign io_VwirePorts_0_14_0_out = Vwire_152_io_out;
  assign io_VwirePorts_0_14_1_out = Vwire_37_io_out;
  assign io_VwirePorts_0_14_3_out = Vwire_129_io_out;
  assign io_VwirePorts_0_14_4_out = Vwire_83_io_out;
  assign io_VwirePorts_0_14_5_out = Vwire_175_io_out;
  assign io_VwirePorts_0_15_0_out = Vwire_153_io_out;
  assign io_VwirePorts_0_15_1_out = Vwire_38_io_out;
  assign io_VwirePorts_0_15_3_out = Vwire_130_io_out;
  assign io_VwirePorts_0_15_4_out = Vwire_84_io_out;
  assign io_VwirePorts_0_15_5_out = Vwire_176_io_out;
  assign io_VwirePorts_0_16_0_out = Vwire_154_io_out;
  assign io_VwirePorts_0_16_1_out = Vwire_39_io_out;
  assign io_VwirePorts_0_16_3_out = Vwire_131_io_out;
  assign io_VwirePorts_0_16_4_out = Vwire_85_io_out;
  assign io_VwirePorts_0_16_5_out = Vwire_177_io_out;
  assign io_VwirePorts_0_17_0_out = Vwire_155_io_out;
  assign io_VwirePorts_0_17_1_out = Vwire_40_io_out;
  assign io_VwirePorts_0_17_3_out = Vwire_132_io_out;
  assign io_VwirePorts_0_17_4_out = Vwire_86_io_out;
  assign io_VwirePorts_0_17_5_out = Vwire_178_io_out;
  assign io_VwirePorts_0_18_0_out = Vwire_156_io_out;
  assign io_VwirePorts_0_18_1_out = Vwire_41_io_out;
  assign io_VwirePorts_0_18_3_out = Vwire_133_io_out;
  assign io_VwirePorts_0_18_4_out = Vwire_87_io_out;
  assign io_VwirePorts_0_18_5_out = Vwire_179_io_out;
  assign io_VwirePorts_0_19_0_out = Vwire_157_io_out;
  assign io_VwirePorts_0_19_1_out = Vwire_42_io_out;
  assign io_VwirePorts_0_19_3_out = Vwire_134_io_out;
  assign io_VwirePorts_0_19_4_out = Vwire_88_io_out;
  assign io_VwirePorts_0_19_5_out = Vwire_180_io_out;
  assign io_VwirePorts_0_20_0_out = Vwire_158_io_out;
  assign io_VwirePorts_0_20_1_out = Vwire_43_io_out;
  assign io_VwirePorts_0_20_3_out = Vwire_135_io_out;
  assign io_VwirePorts_0_20_4_out = Vwire_89_io_out;
  assign io_VwirePorts_0_20_5_out = Vwire_181_io_out;
  assign io_VwirePorts_0_21_0_out = Vwire_159_io_out;
  assign io_VwirePorts_0_21_1_out = Vwire_44_io_out;
  assign io_VwirePorts_0_21_3_out = Vwire_136_io_out;
  assign io_VwirePorts_0_21_4_out = Vwire_90_io_out;
  assign io_VwirePorts_0_21_5_out = Vwire_182_io_out;
  assign io_VwirePorts_0_22_0_out = Vwire_160_io_out;
  assign io_VwirePorts_0_22_1_out = Vwire_45_io_out;
  assign io_VwirePorts_0_22_3_out = Vwire_137_io_out;
  assign io_VwirePorts_0_22_4_out = Vwire_91_io_out;
  assign io_VwirePorts_0_22_5_out = Vwire_183_io_out;
  assign io_VwirePorts_1_0_0_out = Vwire_23_io_out;
  assign io_VwirePorts_1_0_1_out = Vwire_138_io_out;
  assign io_VwirePorts_1_0_2_out = Vwire_92_io_out;
  assign io_VwirePorts_1_0_3_out = Vwire_115_io_out;
  assign io_VwirePorts_1_0_4_out = Vwire_69_io_out;
  assign io_VwirePorts_1_0_5_out = Vwire_161_io_out;
  assign io_VwirePorts_1_1_0_out = Vwire_24_io_out;
  assign io_VwirePorts_1_1_1_out = Vwire_139_io_out;
  assign io_VwirePorts_1_1_2_out = Vwire_93_io_out;
  assign io_VwirePorts_1_1_3_out = Vwire_116_io_out;
  assign io_VwirePorts_1_1_4_out = Vwire_70_io_out;
  assign io_VwirePorts_1_1_5_out = Vwire_162_io_out;
  assign io_VwirePorts_1_2_0_out = Vwire_25_io_out;
  assign io_VwirePorts_1_2_1_out = Vwire_140_io_out;
  assign io_VwirePorts_1_2_2_out = Vwire_94_io_out;
  assign io_VwirePorts_1_2_3_out = Vwire_117_io_out;
  assign io_VwirePorts_1_2_4_out = Vwire_71_io_out;
  assign io_VwirePorts_1_2_5_out = Vwire_163_io_out;
  assign io_VwirePorts_1_3_0_out = Vwire_26_io_out;
  assign io_VwirePorts_1_3_1_out = Vwire_141_io_out;
  assign io_VwirePorts_1_3_2_out = Vwire_95_io_out;
  assign io_VwirePorts_1_3_3_out = Vwire_118_io_out;
  assign io_VwirePorts_1_3_4_out = Vwire_72_io_out;
  assign io_VwirePorts_1_3_5_out = Vwire_164_io_out;
  assign io_VwirePorts_1_4_0_out = Vwire_27_io_out;
  assign io_VwirePorts_1_4_1_out = Vwire_142_io_out;
  assign io_VwirePorts_1_4_2_out = Vwire_96_io_out;
  assign io_VwirePorts_1_4_3_out = Vwire_119_io_out;
  assign io_VwirePorts_1_4_4_out = Vwire_73_io_out;
  assign io_VwirePorts_1_4_5_out = Vwire_165_io_out;
  assign io_VwirePorts_1_5_0_out = Vwire_28_io_out;
  assign io_VwirePorts_1_5_1_out = Vwire_143_io_out;
  assign io_VwirePorts_1_5_2_out = Vwire_97_io_out;
  assign io_VwirePorts_1_5_3_out = Vwire_120_io_out;
  assign io_VwirePorts_1_5_4_out = Vwire_74_io_out;
  assign io_VwirePorts_1_5_5_out = Vwire_166_io_out;
  assign io_VwirePorts_1_6_0_out = Vwire_29_io_out;
  assign io_VwirePorts_1_6_1_out = Vwire_144_io_out;
  assign io_VwirePorts_1_6_2_out = Vwire_98_io_out;
  assign io_VwirePorts_1_6_3_out = Vwire_121_io_out;
  assign io_VwirePorts_1_6_4_out = Vwire_75_io_out;
  assign io_VwirePorts_1_6_5_out = Vwire_167_io_out;
  assign io_VwirePorts_1_7_0_out = Vwire_30_io_out;
  assign io_VwirePorts_1_7_1_out = Vwire_145_io_out;
  assign io_VwirePorts_1_7_2_out = Vwire_99_io_out;
  assign io_VwirePorts_1_7_3_out = Vwire_122_io_out;
  assign io_VwirePorts_1_7_4_out = Vwire_76_io_out;
  assign io_VwirePorts_1_7_5_out = Vwire_168_io_out;
  assign io_VwirePorts_1_8_0_out = Vwire_31_io_out;
  assign io_VwirePorts_1_8_1_out = Vwire_146_io_out;
  assign io_VwirePorts_1_8_2_out = Vwire_100_io_out;
  assign io_VwirePorts_1_8_3_out = Vwire_123_io_out;
  assign io_VwirePorts_1_8_4_out = Vwire_77_io_out;
  assign io_VwirePorts_1_8_5_out = Vwire_169_io_out;
  assign io_VwirePorts_1_9_0_out = Vwire_32_io_out;
  assign io_VwirePorts_1_9_1_out = Vwire_147_io_out;
  assign io_VwirePorts_1_9_2_out = Vwire_101_io_out;
  assign io_VwirePorts_1_9_3_out = Vwire_124_io_out;
  assign io_VwirePorts_1_9_4_out = Vwire_78_io_out;
  assign io_VwirePorts_1_9_5_out = Vwire_170_io_out;
  assign io_VwirePorts_1_10_0_out = Vwire_33_io_out;
  assign io_VwirePorts_1_10_1_out = Vwire_148_io_out;
  assign io_VwirePorts_1_10_2_out = Vwire_102_io_out;
  assign io_VwirePorts_1_10_3_out = Vwire_125_io_out;
  assign io_VwirePorts_1_10_4_out = Vwire_79_io_out;
  assign io_VwirePorts_1_10_5_out = Vwire_171_io_out;
  assign io_VwirePorts_1_11_0_out = Vwire_34_io_out;
  assign io_VwirePorts_1_11_1_out = Vwire_149_io_out;
  assign io_VwirePorts_1_11_2_out = Vwire_103_io_out;
  assign io_VwirePorts_1_11_3_out = Vwire_126_io_out;
  assign io_VwirePorts_1_11_4_out = Vwire_80_io_out;
  assign io_VwirePorts_1_11_5_out = Vwire_172_io_out;
  assign io_VwirePorts_1_12_0_out = Vwire_35_io_out;
  assign io_VwirePorts_1_12_1_out = Vwire_150_io_out;
  assign io_VwirePorts_1_12_2_out = Vwire_104_io_out;
  assign io_VwirePorts_1_12_3_out = Vwire_127_io_out;
  assign io_VwirePorts_1_12_4_out = Vwire_81_io_out;
  assign io_VwirePorts_1_12_5_out = Vwire_173_io_out;
  assign io_VwirePorts_1_13_0_out = Vwire_36_io_out;
  assign io_VwirePorts_1_13_1_out = Vwire_151_io_out;
  assign io_VwirePorts_1_13_2_out = Vwire_105_io_out;
  assign io_VwirePorts_1_13_3_out = Vwire_128_io_out;
  assign io_VwirePorts_1_13_4_out = Vwire_82_io_out;
  assign io_VwirePorts_1_13_5_out = Vwire_174_io_out;
  assign io_VwirePorts_1_14_0_out = Vwire_37_io_out;
  assign io_VwirePorts_1_14_1_out = Vwire_152_io_out;
  assign io_VwirePorts_1_14_2_out = Vwire_106_io_out;
  assign io_VwirePorts_1_14_3_out = Vwire_129_io_out;
  assign io_VwirePorts_1_14_4_out = Vwire_83_io_out;
  assign io_VwirePorts_1_14_5_out = Vwire_175_io_out;
  assign io_VwirePorts_1_15_0_out = Vwire_38_io_out;
  assign io_VwirePorts_1_15_1_out = Vwire_153_io_out;
  assign io_VwirePorts_1_15_2_out = Vwire_107_io_out;
  assign io_VwirePorts_1_15_3_out = Vwire_130_io_out;
  assign io_VwirePorts_1_15_4_out = Vwire_84_io_out;
  assign io_VwirePorts_1_15_5_out = Vwire_176_io_out;
  assign io_VwirePorts_1_16_0_out = Vwire_39_io_out;
  assign io_VwirePorts_1_16_1_out = Vwire_154_io_out;
  assign io_VwirePorts_1_16_2_out = Vwire_108_io_out;
  assign io_VwirePorts_1_16_3_out = Vwire_131_io_out;
  assign io_VwirePorts_1_16_4_out = Vwire_85_io_out;
  assign io_VwirePorts_1_16_5_out = Vwire_177_io_out;
  assign io_VwirePorts_1_17_0_out = Vwire_40_io_out;
  assign io_VwirePorts_1_17_1_out = Vwire_155_io_out;
  assign io_VwirePorts_1_17_2_out = Vwire_109_io_out;
  assign io_VwirePorts_1_17_3_out = Vwire_132_io_out;
  assign io_VwirePorts_1_17_4_out = Vwire_86_io_out;
  assign io_VwirePorts_1_17_5_out = Vwire_178_io_out;
  assign io_VwirePorts_1_18_0_out = Vwire_41_io_out;
  assign io_VwirePorts_1_18_1_out = Vwire_156_io_out;
  assign io_VwirePorts_1_18_2_out = Vwire_110_io_out;
  assign io_VwirePorts_1_18_3_out = Vwire_133_io_out;
  assign io_VwirePorts_1_18_4_out = Vwire_87_io_out;
  assign io_VwirePorts_1_18_5_out = Vwire_179_io_out;
  assign io_VwirePorts_1_19_0_out = Vwire_42_io_out;
  assign io_VwirePorts_1_19_1_out = Vwire_157_io_out;
  assign io_VwirePorts_1_19_2_out = Vwire_111_io_out;
  assign io_VwirePorts_1_19_3_out = Vwire_134_io_out;
  assign io_VwirePorts_1_19_4_out = Vwire_88_io_out;
  assign io_VwirePorts_1_19_5_out = Vwire_180_io_out;
  assign io_VwirePorts_1_20_0_out = Vwire_43_io_out;
  assign io_VwirePorts_1_20_1_out = Vwire_158_io_out;
  assign io_VwirePorts_1_20_2_out = Vwire_112_io_out;
  assign io_VwirePorts_1_20_3_out = Vwire_135_io_out;
  assign io_VwirePorts_1_20_4_out = Vwire_89_io_out;
  assign io_VwirePorts_1_20_5_out = Vwire_181_io_out;
  assign io_VwirePorts_1_21_0_out = Vwire_44_io_out;
  assign io_VwirePorts_1_21_1_out = Vwire_159_io_out;
  assign io_VwirePorts_1_21_2_out = Vwire_113_io_out;
  assign io_VwirePorts_1_21_3_out = Vwire_136_io_out;
  assign io_VwirePorts_1_21_4_out = Vwire_90_io_out;
  assign io_VwirePorts_1_21_5_out = Vwire_182_io_out;
  assign io_VwirePorts_1_22_0_out = Vwire_45_io_out;
  assign io_VwirePorts_1_22_1_out = Vwire_160_io_out;
  assign io_VwirePorts_1_22_2_out = Vwire_114_io_out;
  assign io_VwirePorts_1_22_3_out = Vwire_137_io_out;
  assign io_VwirePorts_1_22_4_out = Vwire_91_io_out;
  assign io_VwirePorts_1_22_5_out = Vwire_183_io_out;
  assign io_VwirePorts_2_0_0_out = Vwire_io_out;
  assign io_VwirePorts_2_0_1_out = Vwire_138_io_out;
  assign io_VwirePorts_2_0_2_out = Vwire_115_io_out;
  assign io_VwirePorts_2_0_3_out = Vwire_92_io_out;
  assign io_VwirePorts_2_0_4_out = Vwire_46_io_out;
  assign io_VwirePorts_2_0_5_out = Vwire_161_io_out;
  assign io_VwirePorts_2_1_0_out = Vwire_1_io_out;
  assign io_VwirePorts_2_1_1_out = Vwire_139_io_out;
  assign io_VwirePorts_2_1_2_out = Vwire_116_io_out;
  assign io_VwirePorts_2_1_3_out = Vwire_93_io_out;
  assign io_VwirePorts_2_1_4_out = Vwire_47_io_out;
  assign io_VwirePorts_2_1_5_out = Vwire_162_io_out;
  assign io_VwirePorts_2_2_0_out = Vwire_2_io_out;
  assign io_VwirePorts_2_2_1_out = Vwire_140_io_out;
  assign io_VwirePorts_2_2_2_out = Vwire_117_io_out;
  assign io_VwirePorts_2_2_3_out = Vwire_94_io_out;
  assign io_VwirePorts_2_2_4_out = Vwire_48_io_out;
  assign io_VwirePorts_2_2_5_out = Vwire_163_io_out;
  assign io_VwirePorts_2_3_0_out = Vwire_3_io_out;
  assign io_VwirePorts_2_3_1_out = Vwire_141_io_out;
  assign io_VwirePorts_2_3_2_out = Vwire_118_io_out;
  assign io_VwirePorts_2_3_3_out = Vwire_95_io_out;
  assign io_VwirePorts_2_3_4_out = Vwire_49_io_out;
  assign io_VwirePorts_2_3_5_out = Vwire_164_io_out;
  assign io_VwirePorts_2_4_0_out = Vwire_4_io_out;
  assign io_VwirePorts_2_4_1_out = Vwire_142_io_out;
  assign io_VwirePorts_2_4_2_out = Vwire_119_io_out;
  assign io_VwirePorts_2_4_3_out = Vwire_96_io_out;
  assign io_VwirePorts_2_4_4_out = Vwire_50_io_out;
  assign io_VwirePorts_2_4_5_out = Vwire_165_io_out;
  assign io_VwirePorts_2_5_0_out = Vwire_5_io_out;
  assign io_VwirePorts_2_5_1_out = Vwire_143_io_out;
  assign io_VwirePorts_2_5_2_out = Vwire_120_io_out;
  assign io_VwirePorts_2_5_3_out = Vwire_97_io_out;
  assign io_VwirePorts_2_5_4_out = Vwire_51_io_out;
  assign io_VwirePorts_2_5_5_out = Vwire_166_io_out;
  assign io_VwirePorts_2_6_0_out = Vwire_6_io_out;
  assign io_VwirePorts_2_6_1_out = Vwire_144_io_out;
  assign io_VwirePorts_2_6_2_out = Vwire_121_io_out;
  assign io_VwirePorts_2_6_3_out = Vwire_98_io_out;
  assign io_VwirePorts_2_6_4_out = Vwire_52_io_out;
  assign io_VwirePorts_2_6_5_out = Vwire_167_io_out;
  assign io_VwirePorts_2_7_0_out = Vwire_7_io_out;
  assign io_VwirePorts_2_7_1_out = Vwire_145_io_out;
  assign io_VwirePorts_2_7_2_out = Vwire_122_io_out;
  assign io_VwirePorts_2_7_3_out = Vwire_99_io_out;
  assign io_VwirePorts_2_7_4_out = Vwire_53_io_out;
  assign io_VwirePorts_2_7_5_out = Vwire_168_io_out;
  assign io_VwirePorts_2_8_0_out = Vwire_8_io_out;
  assign io_VwirePorts_2_8_1_out = Vwire_146_io_out;
  assign io_VwirePorts_2_8_2_out = Vwire_123_io_out;
  assign io_VwirePorts_2_8_3_out = Vwire_100_io_out;
  assign io_VwirePorts_2_8_4_out = Vwire_54_io_out;
  assign io_VwirePorts_2_8_5_out = Vwire_169_io_out;
  assign io_VwirePorts_2_9_0_out = Vwire_9_io_out;
  assign io_VwirePorts_2_9_1_out = Vwire_147_io_out;
  assign io_VwirePorts_2_9_2_out = Vwire_124_io_out;
  assign io_VwirePorts_2_9_3_out = Vwire_101_io_out;
  assign io_VwirePorts_2_9_4_out = Vwire_55_io_out;
  assign io_VwirePorts_2_9_5_out = Vwire_170_io_out;
  assign io_VwirePorts_2_10_0_out = Vwire_10_io_out;
  assign io_VwirePorts_2_10_1_out = Vwire_148_io_out;
  assign io_VwirePorts_2_10_2_out = Vwire_125_io_out;
  assign io_VwirePorts_2_10_3_out = Vwire_102_io_out;
  assign io_VwirePorts_2_10_4_out = Vwire_56_io_out;
  assign io_VwirePorts_2_10_5_out = Vwire_171_io_out;
  assign io_VwirePorts_2_11_0_out = Vwire_11_io_out;
  assign io_VwirePorts_2_11_1_out = Vwire_149_io_out;
  assign io_VwirePorts_2_11_2_out = Vwire_126_io_out;
  assign io_VwirePorts_2_11_3_out = Vwire_103_io_out;
  assign io_VwirePorts_2_11_4_out = Vwire_57_io_out;
  assign io_VwirePorts_2_11_5_out = Vwire_172_io_out;
  assign io_VwirePorts_2_12_0_out = Vwire_12_io_out;
  assign io_VwirePorts_2_12_1_out = Vwire_150_io_out;
  assign io_VwirePorts_2_12_2_out = Vwire_127_io_out;
  assign io_VwirePorts_2_12_3_out = Vwire_104_io_out;
  assign io_VwirePorts_2_12_4_out = Vwire_58_io_out;
  assign io_VwirePorts_2_12_5_out = Vwire_173_io_out;
  assign io_VwirePorts_2_13_0_out = Vwire_13_io_out;
  assign io_VwirePorts_2_13_1_out = Vwire_151_io_out;
  assign io_VwirePorts_2_13_2_out = Vwire_128_io_out;
  assign io_VwirePorts_2_13_3_out = Vwire_105_io_out;
  assign io_VwirePorts_2_13_4_out = Vwire_59_io_out;
  assign io_VwirePorts_2_13_5_out = Vwire_174_io_out;
  assign io_VwirePorts_2_14_0_out = Vwire_14_io_out;
  assign io_VwirePorts_2_14_1_out = Vwire_152_io_out;
  assign io_VwirePorts_2_14_2_out = Vwire_129_io_out;
  assign io_VwirePorts_2_14_3_out = Vwire_106_io_out;
  assign io_VwirePorts_2_14_4_out = Vwire_60_io_out;
  assign io_VwirePorts_2_14_5_out = Vwire_175_io_out;
  assign io_VwirePorts_2_15_0_out = Vwire_15_io_out;
  assign io_VwirePorts_2_15_1_out = Vwire_153_io_out;
  assign io_VwirePorts_2_15_2_out = Vwire_130_io_out;
  assign io_VwirePorts_2_15_3_out = Vwire_107_io_out;
  assign io_VwirePorts_2_15_4_out = Vwire_61_io_out;
  assign io_VwirePorts_2_15_5_out = Vwire_176_io_out;
  assign io_VwirePorts_2_16_0_out = Vwire_16_io_out;
  assign io_VwirePorts_2_16_1_out = Vwire_154_io_out;
  assign io_VwirePorts_2_16_2_out = Vwire_131_io_out;
  assign io_VwirePorts_2_16_3_out = Vwire_108_io_out;
  assign io_VwirePorts_2_16_4_out = Vwire_62_io_out;
  assign io_VwirePorts_2_16_5_out = Vwire_177_io_out;
  assign io_VwirePorts_2_17_0_out = Vwire_17_io_out;
  assign io_VwirePorts_2_17_1_out = Vwire_155_io_out;
  assign io_VwirePorts_2_17_2_out = Vwire_132_io_out;
  assign io_VwirePorts_2_17_3_out = Vwire_109_io_out;
  assign io_VwirePorts_2_17_4_out = Vwire_63_io_out;
  assign io_VwirePorts_2_17_5_out = Vwire_178_io_out;
  assign io_VwirePorts_2_18_0_out = Vwire_18_io_out;
  assign io_VwirePorts_2_18_1_out = Vwire_156_io_out;
  assign io_VwirePorts_2_18_2_out = Vwire_133_io_out;
  assign io_VwirePorts_2_18_3_out = Vwire_110_io_out;
  assign io_VwirePorts_2_18_4_out = Vwire_64_io_out;
  assign io_VwirePorts_2_18_5_out = Vwire_179_io_out;
  assign io_VwirePorts_2_19_0_out = Vwire_19_io_out;
  assign io_VwirePorts_2_19_1_out = Vwire_157_io_out;
  assign io_VwirePorts_2_19_2_out = Vwire_134_io_out;
  assign io_VwirePorts_2_19_3_out = Vwire_111_io_out;
  assign io_VwirePorts_2_19_4_out = Vwire_65_io_out;
  assign io_VwirePorts_2_19_5_out = Vwire_180_io_out;
  assign io_VwirePorts_2_20_0_out = Vwire_20_io_out;
  assign io_VwirePorts_2_20_1_out = Vwire_158_io_out;
  assign io_VwirePorts_2_20_2_out = Vwire_135_io_out;
  assign io_VwirePorts_2_20_3_out = Vwire_112_io_out;
  assign io_VwirePorts_2_20_4_out = Vwire_66_io_out;
  assign io_VwirePorts_2_20_5_out = Vwire_181_io_out;
  assign io_VwirePorts_2_21_0_out = Vwire_21_io_out;
  assign io_VwirePorts_2_21_1_out = Vwire_159_io_out;
  assign io_VwirePorts_2_21_2_out = Vwire_136_io_out;
  assign io_VwirePorts_2_21_3_out = Vwire_113_io_out;
  assign io_VwirePorts_2_21_4_out = Vwire_67_io_out;
  assign io_VwirePorts_2_21_5_out = Vwire_182_io_out;
  assign io_VwirePorts_2_22_0_out = Vwire_22_io_out;
  assign io_VwirePorts_2_22_1_out = Vwire_160_io_out;
  assign io_VwirePorts_2_22_2_out = Vwire_137_io_out;
  assign io_VwirePorts_2_22_3_out = Vwire_114_io_out;
  assign io_VwirePorts_2_22_4_out = Vwire_68_io_out;
  assign io_VwirePorts_2_22_5_out = Vwire_183_io_out;
  assign io_VwirePorts_3_0_0_out = Vwire_138_io_out;
  assign io_VwirePorts_3_0_1_out = Vwire_io_out;
  assign io_VwirePorts_3_0_3_out = Vwire_92_io_out;
  assign io_VwirePorts_3_0_4_out = Vwire_46_io_out;
  assign io_VwirePorts_3_0_5_out = Vwire_161_io_out;
  assign io_VwirePorts_3_1_0_out = Vwire_139_io_out;
  assign io_VwirePorts_3_1_1_out = Vwire_1_io_out;
  assign io_VwirePorts_3_1_3_out = Vwire_93_io_out;
  assign io_VwirePorts_3_1_4_out = Vwire_47_io_out;
  assign io_VwirePorts_3_1_5_out = Vwire_162_io_out;
  assign io_VwirePorts_3_2_0_out = Vwire_140_io_out;
  assign io_VwirePorts_3_2_1_out = Vwire_2_io_out;
  assign io_VwirePorts_3_2_3_out = Vwire_94_io_out;
  assign io_VwirePorts_3_2_4_out = Vwire_48_io_out;
  assign io_VwirePorts_3_2_5_out = Vwire_163_io_out;
  assign io_VwirePorts_3_3_0_out = Vwire_141_io_out;
  assign io_VwirePorts_3_3_1_out = Vwire_3_io_out;
  assign io_VwirePorts_3_3_3_out = Vwire_95_io_out;
  assign io_VwirePorts_3_3_4_out = Vwire_49_io_out;
  assign io_VwirePorts_3_3_5_out = Vwire_164_io_out;
  assign io_VwirePorts_3_4_0_out = Vwire_142_io_out;
  assign io_VwirePorts_3_4_1_out = Vwire_4_io_out;
  assign io_VwirePorts_3_4_3_out = Vwire_96_io_out;
  assign io_VwirePorts_3_4_4_out = Vwire_50_io_out;
  assign io_VwirePorts_3_4_5_out = Vwire_165_io_out;
  assign io_VwirePorts_3_5_0_out = Vwire_143_io_out;
  assign io_VwirePorts_3_5_1_out = Vwire_5_io_out;
  assign io_VwirePorts_3_5_3_out = Vwire_97_io_out;
  assign io_VwirePorts_3_5_4_out = Vwire_51_io_out;
  assign io_VwirePorts_3_5_5_out = Vwire_166_io_out;
  assign io_VwirePorts_3_6_0_out = Vwire_144_io_out;
  assign io_VwirePorts_3_6_1_out = Vwire_6_io_out;
  assign io_VwirePorts_3_6_3_out = Vwire_98_io_out;
  assign io_VwirePorts_3_6_4_out = Vwire_52_io_out;
  assign io_VwirePorts_3_6_5_out = Vwire_167_io_out;
  assign io_VwirePorts_3_7_0_out = Vwire_145_io_out;
  assign io_VwirePorts_3_7_1_out = Vwire_7_io_out;
  assign io_VwirePorts_3_7_3_out = Vwire_99_io_out;
  assign io_VwirePorts_3_7_4_out = Vwire_53_io_out;
  assign io_VwirePorts_3_7_5_out = Vwire_168_io_out;
  assign io_VwirePorts_3_8_0_out = Vwire_146_io_out;
  assign io_VwirePorts_3_8_1_out = Vwire_8_io_out;
  assign io_VwirePorts_3_8_3_out = Vwire_100_io_out;
  assign io_VwirePorts_3_8_4_out = Vwire_54_io_out;
  assign io_VwirePorts_3_8_5_out = Vwire_169_io_out;
  assign io_VwirePorts_3_9_0_out = Vwire_147_io_out;
  assign io_VwirePorts_3_9_1_out = Vwire_9_io_out;
  assign io_VwirePorts_3_9_3_out = Vwire_101_io_out;
  assign io_VwirePorts_3_9_4_out = Vwire_55_io_out;
  assign io_VwirePorts_3_9_5_out = Vwire_170_io_out;
  assign io_VwirePorts_3_10_0_out = Vwire_148_io_out;
  assign io_VwirePorts_3_10_1_out = Vwire_10_io_out;
  assign io_VwirePorts_3_10_3_out = Vwire_102_io_out;
  assign io_VwirePorts_3_10_4_out = Vwire_56_io_out;
  assign io_VwirePorts_3_10_5_out = Vwire_171_io_out;
  assign io_VwirePorts_3_11_0_out = Vwire_149_io_out;
  assign io_VwirePorts_3_11_1_out = Vwire_11_io_out;
  assign io_VwirePorts_3_11_3_out = Vwire_103_io_out;
  assign io_VwirePorts_3_11_4_out = Vwire_57_io_out;
  assign io_VwirePorts_3_11_5_out = Vwire_172_io_out;
  assign io_VwirePorts_3_12_0_out = Vwire_150_io_out;
  assign io_VwirePorts_3_12_1_out = Vwire_12_io_out;
  assign io_VwirePorts_3_12_3_out = Vwire_104_io_out;
  assign io_VwirePorts_3_12_4_out = Vwire_58_io_out;
  assign io_VwirePorts_3_12_5_out = Vwire_173_io_out;
  assign io_VwirePorts_3_13_0_out = Vwire_151_io_out;
  assign io_VwirePorts_3_13_1_out = Vwire_13_io_out;
  assign io_VwirePorts_3_13_3_out = Vwire_105_io_out;
  assign io_VwirePorts_3_13_4_out = Vwire_59_io_out;
  assign io_VwirePorts_3_13_5_out = Vwire_174_io_out;
  assign io_VwirePorts_3_14_0_out = Vwire_152_io_out;
  assign io_VwirePorts_3_14_1_out = Vwire_14_io_out;
  assign io_VwirePorts_3_14_3_out = Vwire_106_io_out;
  assign io_VwirePorts_3_14_4_out = Vwire_60_io_out;
  assign io_VwirePorts_3_14_5_out = Vwire_175_io_out;
  assign io_VwirePorts_3_15_0_out = Vwire_153_io_out;
  assign io_VwirePorts_3_15_1_out = Vwire_15_io_out;
  assign io_VwirePorts_3_15_3_out = Vwire_107_io_out;
  assign io_VwirePorts_3_15_4_out = Vwire_61_io_out;
  assign io_VwirePorts_3_15_5_out = Vwire_176_io_out;
  assign io_VwirePorts_3_16_0_out = Vwire_154_io_out;
  assign io_VwirePorts_3_16_1_out = Vwire_16_io_out;
  assign io_VwirePorts_3_16_3_out = Vwire_108_io_out;
  assign io_VwirePorts_3_16_4_out = Vwire_62_io_out;
  assign io_VwirePorts_3_16_5_out = Vwire_177_io_out;
  assign io_VwirePorts_3_17_0_out = Vwire_155_io_out;
  assign io_VwirePorts_3_17_1_out = Vwire_17_io_out;
  assign io_VwirePorts_3_17_3_out = Vwire_109_io_out;
  assign io_VwirePorts_3_17_4_out = Vwire_63_io_out;
  assign io_VwirePorts_3_17_5_out = Vwire_178_io_out;
  assign io_VwirePorts_3_18_0_out = Vwire_156_io_out;
  assign io_VwirePorts_3_18_1_out = Vwire_18_io_out;
  assign io_VwirePorts_3_18_3_out = Vwire_110_io_out;
  assign io_VwirePorts_3_18_4_out = Vwire_64_io_out;
  assign io_VwirePorts_3_18_5_out = Vwire_179_io_out;
  assign io_VwirePorts_3_19_0_out = Vwire_157_io_out;
  assign io_VwirePorts_3_19_1_out = Vwire_19_io_out;
  assign io_VwirePorts_3_19_3_out = Vwire_111_io_out;
  assign io_VwirePorts_3_19_4_out = Vwire_65_io_out;
  assign io_VwirePorts_3_19_5_out = Vwire_180_io_out;
  assign io_VwirePorts_3_20_0_out = Vwire_158_io_out;
  assign io_VwirePorts_3_20_1_out = Vwire_20_io_out;
  assign io_VwirePorts_3_20_3_out = Vwire_112_io_out;
  assign io_VwirePorts_3_20_4_out = Vwire_66_io_out;
  assign io_VwirePorts_3_20_5_out = Vwire_181_io_out;
  assign io_VwirePorts_3_21_0_out = Vwire_159_io_out;
  assign io_VwirePorts_3_21_1_out = Vwire_21_io_out;
  assign io_VwirePorts_3_21_3_out = Vwire_113_io_out;
  assign io_VwirePorts_3_21_4_out = Vwire_67_io_out;
  assign io_VwirePorts_3_21_5_out = Vwire_182_io_out;
  assign io_VwirePorts_3_22_0_out = Vwire_160_io_out;
  assign io_VwirePorts_3_22_1_out = Vwire_22_io_out;
  assign io_VwirePorts_3_22_3_out = Vwire_114_io_out;
  assign io_VwirePorts_3_22_4_out = Vwire_68_io_out;
  assign io_VwirePorts_3_22_5_out = Vwire_183_io_out;
  Vwire_0 Vwire(
       .io_in_1( io_VwirePorts_3_0_1_in ),
       .io_in_0( io_VwirePorts_2_0_0_in ),
       .io_en_1( io_VwirePorts_3_0_1_en ),
       .io_en_0( io_VwirePorts_2_0_0_en ),
       .io_out( Vwire_io_out )
  );
  Vwire_0 Vwire_1(
       .io_in_1( io_VwirePorts_3_1_1_in ),
       .io_in_0( io_VwirePorts_2_1_0_in ),
       .io_en_1( io_VwirePorts_3_1_1_en ),
       .io_en_0( io_VwirePorts_2_1_0_en ),
       .io_out( Vwire_1_io_out )
  );
  Vwire_0 Vwire_2(
       .io_in_1( io_VwirePorts_3_2_1_in ),
       .io_in_0( io_VwirePorts_2_2_0_in ),
       .io_en_1( io_VwirePorts_3_2_1_en ),
       .io_en_0( io_VwirePorts_2_2_0_en ),
       .io_out( Vwire_2_io_out )
  );
  Vwire_0 Vwire_3(
       .io_in_1( io_VwirePorts_3_3_1_in ),
       .io_in_0( io_VwirePorts_2_3_0_in ),
       .io_en_1( io_VwirePorts_3_3_1_en ),
       .io_en_0( io_VwirePorts_2_3_0_en ),
       .io_out( Vwire_3_io_out )
  );
  Vwire_0 Vwire_4(
       .io_in_1( io_VwirePorts_3_4_1_in ),
       .io_in_0( io_VwirePorts_2_4_0_in ),
       .io_en_1( io_VwirePorts_3_4_1_en ),
       .io_en_0( io_VwirePorts_2_4_0_en ),
       .io_out( Vwire_4_io_out )
  );
  Vwire_0 Vwire_5(
       .io_in_1( io_VwirePorts_3_5_1_in ),
       .io_in_0( io_VwirePorts_2_5_0_in ),
       .io_en_1( io_VwirePorts_3_5_1_en ),
       .io_en_0( io_VwirePorts_2_5_0_en ),
       .io_out( Vwire_5_io_out )
  );
  Vwire_0 Vwire_6(
       .io_in_1( io_VwirePorts_3_6_1_in ),
       .io_in_0( io_VwirePorts_2_6_0_in ),
       .io_en_1( io_VwirePorts_3_6_1_en ),
       .io_en_0( io_VwirePorts_2_6_0_en ),
       .io_out( Vwire_6_io_out )
  );
  Vwire_0 Vwire_7(
       .io_in_1( io_VwirePorts_3_7_1_in ),
       .io_in_0( io_VwirePorts_2_7_0_in ),
       .io_en_1( io_VwirePorts_3_7_1_en ),
       .io_en_0( io_VwirePorts_2_7_0_en ),
       .io_out( Vwire_7_io_out )
  );
  Vwire_0 Vwire_8(
       .io_in_1( io_VwirePorts_3_8_1_in ),
       .io_in_0( io_VwirePorts_2_8_0_in ),
       .io_en_1( io_VwirePorts_3_8_1_en ),
       .io_en_0( io_VwirePorts_2_8_0_en ),
       .io_out( Vwire_8_io_out )
  );
  Vwire_0 Vwire_9(
       .io_in_1( io_VwirePorts_3_9_1_in ),
       .io_in_0( io_VwirePorts_2_9_0_in ),
       .io_en_1( io_VwirePorts_3_9_1_en ),
       .io_en_0( io_VwirePorts_2_9_0_en ),
       .io_out( Vwire_9_io_out )
  );
  Vwire_0 Vwire_10(
       .io_in_1( io_VwirePorts_3_10_1_in ),
       .io_in_0( io_VwirePorts_2_10_0_in ),
       .io_en_1( io_VwirePorts_3_10_1_en ),
       .io_en_0( io_VwirePorts_2_10_0_en ),
       .io_out( Vwire_10_io_out )
  );
  Vwire_0 Vwire_11(
       .io_in_1( io_VwirePorts_3_11_1_in ),
       .io_in_0( io_VwirePorts_2_11_0_in ),
       .io_en_1( io_VwirePorts_3_11_1_en ),
       .io_en_0( io_VwirePorts_2_11_0_en ),
       .io_out( Vwire_11_io_out )
  );
  Vwire_0 Vwire_12(
       .io_in_1( io_VwirePorts_3_12_1_in ),
       .io_in_0( io_VwirePorts_2_12_0_in ),
       .io_en_1( io_VwirePorts_3_12_1_en ),
       .io_en_0( io_VwirePorts_2_12_0_en ),
       .io_out( Vwire_12_io_out )
  );
  Vwire_0 Vwire_13(
       .io_in_1( io_VwirePorts_3_13_1_in ),
       .io_in_0( io_VwirePorts_2_13_0_in ),
       .io_en_1( io_VwirePorts_3_13_1_en ),
       .io_en_0( io_VwirePorts_2_13_0_en ),
       .io_out( Vwire_13_io_out )
  );
  Vwire_0 Vwire_14(
       .io_in_1( io_VwirePorts_3_14_1_in ),
       .io_in_0( io_VwirePorts_2_14_0_in ),
       .io_en_1( io_VwirePorts_3_14_1_en ),
       .io_en_0( io_VwirePorts_2_14_0_en ),
       .io_out( Vwire_14_io_out )
  );
  Vwire_0 Vwire_15(
       .io_in_1( io_VwirePorts_3_15_1_in ),
       .io_in_0( io_VwirePorts_2_15_0_in ),
       .io_en_1( io_VwirePorts_3_15_1_en ),
       .io_en_0( io_VwirePorts_2_15_0_en ),
       .io_out( Vwire_15_io_out )
  );
  Vwire_0 Vwire_16(
       .io_in_1( io_VwirePorts_3_16_1_in ),
       .io_in_0( io_VwirePorts_2_16_0_in ),
       .io_en_1( io_VwirePorts_3_16_1_en ),
       .io_en_0( io_VwirePorts_2_16_0_en ),
       .io_out( Vwire_16_io_out )
  );
  Vwire_0 Vwire_17(
       .io_in_1( io_VwirePorts_3_17_1_in ),
       .io_in_0( io_VwirePorts_2_17_0_in ),
       .io_en_1( io_VwirePorts_3_17_1_en ),
       .io_en_0( io_VwirePorts_2_17_0_en ),
       .io_out( Vwire_17_io_out )
  );
  Vwire_0 Vwire_18(
       .io_in_1( io_VwirePorts_3_18_1_in ),
       .io_in_0( io_VwirePorts_2_18_0_in ),
       .io_en_1( io_VwirePorts_3_18_1_en ),
       .io_en_0( io_VwirePorts_2_18_0_en ),
       .io_out( Vwire_18_io_out )
  );
  Vwire_0 Vwire_19(
       .io_in_1( io_VwirePorts_3_19_1_in ),
       .io_in_0( io_VwirePorts_2_19_0_in ),
       .io_en_1( io_VwirePorts_3_19_1_en ),
       .io_en_0( io_VwirePorts_2_19_0_en ),
       .io_out( Vwire_19_io_out )
  );
  Vwire_0 Vwire_20(
       .io_in_1( io_VwirePorts_3_20_1_in ),
       .io_in_0( io_VwirePorts_2_20_0_in ),
       .io_en_1( io_VwirePorts_3_20_1_en ),
       .io_en_0( io_VwirePorts_2_20_0_en ),
       .io_out( Vwire_20_io_out )
  );
  Vwire_0 Vwire_21(
       .io_in_1( io_VwirePorts_3_21_1_in ),
       .io_in_0( io_VwirePorts_2_21_0_in ),
       .io_en_1( io_VwirePorts_3_21_1_en ),
       .io_en_0( io_VwirePorts_2_21_0_en ),
       .io_out( Vwire_21_io_out )
  );
  Vwire_0 Vwire_22(
       .io_in_1( io_VwirePorts_3_22_1_in ),
       .io_in_0( io_VwirePorts_2_22_0_in ),
       .io_en_1( io_VwirePorts_3_22_1_en ),
       .io_en_0( io_VwirePorts_2_22_0_en ),
       .io_out( Vwire_22_io_out )
  );
  Vwire_0 Vwire_23(
       .io_in_1( io_VwirePorts_1_0_0_in ),
       .io_in_0( io_VwirePorts_0_0_1_in ),
       .io_en_1( io_VwirePorts_1_0_0_en ),
       .io_en_0( io_VwirePorts_0_0_1_en ),
       .io_out( Vwire_23_io_out )
  );
  Vwire_0 Vwire_24(
       .io_in_1( io_VwirePorts_1_1_0_in ),
       .io_in_0( io_VwirePorts_0_1_1_in ),
       .io_en_1( io_VwirePorts_1_1_0_en ),
       .io_en_0( io_VwirePorts_0_1_1_en ),
       .io_out( Vwire_24_io_out )
  );
  Vwire_0 Vwire_25(
       .io_in_1( io_VwirePorts_1_2_0_in ),
       .io_in_0( io_VwirePorts_0_2_1_in ),
       .io_en_1( io_VwirePorts_1_2_0_en ),
       .io_en_0( io_VwirePorts_0_2_1_en ),
       .io_out( Vwire_25_io_out )
  );
  Vwire_0 Vwire_26(
       .io_in_1( io_VwirePorts_1_3_0_in ),
       .io_in_0( io_VwirePorts_0_3_1_in ),
       .io_en_1( io_VwirePorts_1_3_0_en ),
       .io_en_0( io_VwirePorts_0_3_1_en ),
       .io_out( Vwire_26_io_out )
  );
  Vwire_0 Vwire_27(
       .io_in_1( io_VwirePorts_1_4_0_in ),
       .io_in_0( io_VwirePorts_0_4_1_in ),
       .io_en_1( io_VwirePorts_1_4_0_en ),
       .io_en_0( io_VwirePorts_0_4_1_en ),
       .io_out( Vwire_27_io_out )
  );
  Vwire_0 Vwire_28(
       .io_in_1( io_VwirePorts_1_5_0_in ),
       .io_in_0( io_VwirePorts_0_5_1_in ),
       .io_en_1( io_VwirePorts_1_5_0_en ),
       .io_en_0( io_VwirePorts_0_5_1_en ),
       .io_out( Vwire_28_io_out )
  );
  Vwire_0 Vwire_29(
       .io_in_1( io_VwirePorts_1_6_0_in ),
       .io_in_0( io_VwirePorts_0_6_1_in ),
       .io_en_1( io_VwirePorts_1_6_0_en ),
       .io_en_0( io_VwirePorts_0_6_1_en ),
       .io_out( Vwire_29_io_out )
  );
  Vwire_0 Vwire_30(
       .io_in_1( io_VwirePorts_1_7_0_in ),
       .io_in_0( io_VwirePorts_0_7_1_in ),
       .io_en_1( io_VwirePorts_1_7_0_en ),
       .io_en_0( io_VwirePorts_0_7_1_en ),
       .io_out( Vwire_30_io_out )
  );
  Vwire_0 Vwire_31(
       .io_in_1( io_VwirePorts_1_8_0_in ),
       .io_in_0( io_VwirePorts_0_8_1_in ),
       .io_en_1( io_VwirePorts_1_8_0_en ),
       .io_en_0( io_VwirePorts_0_8_1_en ),
       .io_out( Vwire_31_io_out )
  );
  Vwire_0 Vwire_32(
       .io_in_1( io_VwirePorts_1_9_0_in ),
       .io_in_0( io_VwirePorts_0_9_1_in ),
       .io_en_1( io_VwirePorts_1_9_0_en ),
       .io_en_0( io_VwirePorts_0_9_1_en ),
       .io_out( Vwire_32_io_out )
  );
  Vwire_0 Vwire_33(
       .io_in_1( io_VwirePorts_1_10_0_in ),
       .io_in_0( io_VwirePorts_0_10_1_in ),
       .io_en_1( io_VwirePorts_1_10_0_en ),
       .io_en_0( io_VwirePorts_0_10_1_en ),
       .io_out( Vwire_33_io_out )
  );
  Vwire_0 Vwire_34(
       .io_in_1( io_VwirePorts_1_11_0_in ),
       .io_in_0( io_VwirePorts_0_11_1_in ),
       .io_en_1( io_VwirePorts_1_11_0_en ),
       .io_en_0( io_VwirePorts_0_11_1_en ),
       .io_out( Vwire_34_io_out )
  );
  Vwire_0 Vwire_35(
       .io_in_1( io_VwirePorts_1_12_0_in ),
       .io_in_0( io_VwirePorts_0_12_1_in ),
       .io_en_1( io_VwirePorts_1_12_0_en ),
       .io_en_0( io_VwirePorts_0_12_1_en ),
       .io_out( Vwire_35_io_out )
  );
  Vwire_0 Vwire_36(
       .io_in_1( io_VwirePorts_1_13_0_in ),
       .io_in_0( io_VwirePorts_0_13_1_in ),
       .io_en_1( io_VwirePorts_1_13_0_en ),
       .io_en_0( io_VwirePorts_0_13_1_en ),
       .io_out( Vwire_36_io_out )
  );
  Vwire_0 Vwire_37(
       .io_in_1( io_VwirePorts_1_14_0_in ),
       .io_in_0( io_VwirePorts_0_14_1_in ),
       .io_en_1( io_VwirePorts_1_14_0_en ),
       .io_en_0( io_VwirePorts_0_14_1_en ),
       .io_out( Vwire_37_io_out )
  );
  Vwire_0 Vwire_38(
       .io_in_1( io_VwirePorts_1_15_0_in ),
       .io_in_0( io_VwirePorts_0_15_1_in ),
       .io_en_1( io_VwirePorts_1_15_0_en ),
       .io_en_0( io_VwirePorts_0_15_1_en ),
       .io_out( Vwire_38_io_out )
  );
  Vwire_0 Vwire_39(
       .io_in_1( io_VwirePorts_1_16_0_in ),
       .io_in_0( io_VwirePorts_0_16_1_in ),
       .io_en_1( io_VwirePorts_1_16_0_en ),
       .io_en_0( io_VwirePorts_0_16_1_en ),
       .io_out( Vwire_39_io_out )
  );
  Vwire_0 Vwire_40(
       .io_in_1( io_VwirePorts_1_17_0_in ),
       .io_in_0( io_VwirePorts_0_17_1_in ),
       .io_en_1( io_VwirePorts_1_17_0_en ),
       .io_en_0( io_VwirePorts_0_17_1_en ),
       .io_out( Vwire_40_io_out )
  );
  Vwire_0 Vwire_41(
       .io_in_1( io_VwirePorts_1_18_0_in ),
       .io_in_0( io_VwirePorts_0_18_1_in ),
       .io_en_1( io_VwirePorts_1_18_0_en ),
       .io_en_0( io_VwirePorts_0_18_1_en ),
       .io_out( Vwire_41_io_out )
  );
  Vwire_0 Vwire_42(
       .io_in_1( io_VwirePorts_1_19_0_in ),
       .io_in_0( io_VwirePorts_0_19_1_in ),
       .io_en_1( io_VwirePorts_1_19_0_en ),
       .io_en_0( io_VwirePorts_0_19_1_en ),
       .io_out( Vwire_42_io_out )
  );
  Vwire_0 Vwire_43(
       .io_in_1( io_VwirePorts_1_20_0_in ),
       .io_in_0( io_VwirePorts_0_20_1_in ),
       .io_en_1( io_VwirePorts_1_20_0_en ),
       .io_en_0( io_VwirePorts_0_20_1_en ),
       .io_out( Vwire_43_io_out )
  );
  Vwire_0 Vwire_44(
       .io_in_1( io_VwirePorts_1_21_0_in ),
       .io_in_0( io_VwirePorts_0_21_1_in ),
       .io_en_1( io_VwirePorts_1_21_0_en ),
       .io_en_0( io_VwirePorts_0_21_1_en ),
       .io_out( Vwire_44_io_out )
  );
  Vwire_0 Vwire_45(
       .io_in_1( io_VwirePorts_1_22_0_in ),
       .io_in_0( io_VwirePorts_0_22_1_in ),
       .io_en_1( io_VwirePorts_1_22_0_en ),
       .io_en_0( io_VwirePorts_0_22_1_en ),
       .io_out( Vwire_45_io_out )
  );
  Vwire_0 Vwire_46(
       .io_in_1( io_VwirePorts_3_0_4_in ),
       .io_in_0( io_VwirePorts_2_0_4_in ),
       .io_en_1( io_VwirePorts_3_0_4_en ),
       .io_en_0( io_VwirePorts_2_0_4_en ),
       .io_out( Vwire_46_io_out )
  );
  Vwire_0 Vwire_47(
       .io_in_1( io_VwirePorts_3_1_4_in ),
       .io_in_0( io_VwirePorts_2_1_4_in ),
       .io_en_1( io_VwirePorts_3_1_4_en ),
       .io_en_0( io_VwirePorts_2_1_4_en ),
       .io_out( Vwire_47_io_out )
  );
  Vwire_0 Vwire_48(
       .io_in_1( io_VwirePorts_3_2_4_in ),
       .io_in_0( io_VwirePorts_2_2_4_in ),
       .io_en_1( io_VwirePorts_3_2_4_en ),
       .io_en_0( io_VwirePorts_2_2_4_en ),
       .io_out( Vwire_48_io_out )
  );
  Vwire_0 Vwire_49(
       .io_in_1( io_VwirePorts_3_3_4_in ),
       .io_in_0( io_VwirePorts_2_3_4_in ),
       .io_en_1( io_VwirePorts_3_3_4_en ),
       .io_en_0( io_VwirePorts_2_3_4_en ),
       .io_out( Vwire_49_io_out )
  );
  Vwire_0 Vwire_50(
       .io_in_1( io_VwirePorts_3_4_4_in ),
       .io_in_0( io_VwirePorts_2_4_4_in ),
       .io_en_1( io_VwirePorts_3_4_4_en ),
       .io_en_0( io_VwirePorts_2_4_4_en ),
       .io_out( Vwire_50_io_out )
  );
  Vwire_0 Vwire_51(
       .io_in_1( io_VwirePorts_3_5_4_in ),
       .io_in_0( io_VwirePorts_2_5_4_in ),
       .io_en_1( io_VwirePorts_3_5_4_en ),
       .io_en_0( io_VwirePorts_2_5_4_en ),
       .io_out( Vwire_51_io_out )
  );
  Vwire_0 Vwire_52(
       .io_in_1( io_VwirePorts_3_6_4_in ),
       .io_in_0( io_VwirePorts_2_6_4_in ),
       .io_en_1( io_VwirePorts_3_6_4_en ),
       .io_en_0( io_VwirePorts_2_6_4_en ),
       .io_out( Vwire_52_io_out )
  );
  Vwire_0 Vwire_53(
       .io_in_1( io_VwirePorts_3_7_4_in ),
       .io_in_0( io_VwirePorts_2_7_4_in ),
       .io_en_1( io_VwirePorts_3_7_4_en ),
       .io_en_0( io_VwirePorts_2_7_4_en ),
       .io_out( Vwire_53_io_out )
  );
  Vwire_0 Vwire_54(
       .io_in_1( io_VwirePorts_3_8_4_in ),
       .io_in_0( io_VwirePorts_2_8_4_in ),
       .io_en_1( io_VwirePorts_3_8_4_en ),
       .io_en_0( io_VwirePorts_2_8_4_en ),
       .io_out( Vwire_54_io_out )
  );
  Vwire_0 Vwire_55(
       .io_in_1( io_VwirePorts_3_9_4_in ),
       .io_in_0( io_VwirePorts_2_9_4_in ),
       .io_en_1( io_VwirePorts_3_9_4_en ),
       .io_en_0( io_VwirePorts_2_9_4_en ),
       .io_out( Vwire_55_io_out )
  );
  Vwire_0 Vwire_56(
       .io_in_1( io_VwirePorts_3_10_4_in ),
       .io_in_0( io_VwirePorts_2_10_4_in ),
       .io_en_1( io_VwirePorts_3_10_4_en ),
       .io_en_0( io_VwirePorts_2_10_4_en ),
       .io_out( Vwire_56_io_out )
  );
  Vwire_0 Vwire_57(
       .io_in_1( io_VwirePorts_3_11_4_in ),
       .io_in_0( io_VwirePorts_2_11_4_in ),
       .io_en_1( io_VwirePorts_3_11_4_en ),
       .io_en_0( io_VwirePorts_2_11_4_en ),
       .io_out( Vwire_57_io_out )
  );
  Vwire_0 Vwire_58(
       .io_in_1( io_VwirePorts_3_12_4_in ),
       .io_in_0( io_VwirePorts_2_12_4_in ),
       .io_en_1( io_VwirePorts_3_12_4_en ),
       .io_en_0( io_VwirePorts_2_12_4_en ),
       .io_out( Vwire_58_io_out )
  );
  Vwire_0 Vwire_59(
       .io_in_1( io_VwirePorts_3_13_4_in ),
       .io_in_0( io_VwirePorts_2_13_4_in ),
       .io_en_1( io_VwirePorts_3_13_4_en ),
       .io_en_0( io_VwirePorts_2_13_4_en ),
       .io_out( Vwire_59_io_out )
  );
  Vwire_0 Vwire_60(
       .io_in_1( io_VwirePorts_3_14_4_in ),
       .io_in_0( io_VwirePorts_2_14_4_in ),
       .io_en_1( io_VwirePorts_3_14_4_en ),
       .io_en_0( io_VwirePorts_2_14_4_en ),
       .io_out( Vwire_60_io_out )
  );
  Vwire_0 Vwire_61(
       .io_in_1( io_VwirePorts_3_15_4_in ),
       .io_in_0( io_VwirePorts_2_15_4_in ),
       .io_en_1( io_VwirePorts_3_15_4_en ),
       .io_en_0( io_VwirePorts_2_15_4_en ),
       .io_out( Vwire_61_io_out )
  );
  Vwire_0 Vwire_62(
       .io_in_1( io_VwirePorts_3_16_4_in ),
       .io_in_0( io_VwirePorts_2_16_4_in ),
       .io_en_1( io_VwirePorts_3_16_4_en ),
       .io_en_0( io_VwirePorts_2_16_4_en ),
       .io_out( Vwire_62_io_out )
  );
  Vwire_0 Vwire_63(
       .io_in_1( io_VwirePorts_3_17_4_in ),
       .io_in_0( io_VwirePorts_2_17_4_in ),
       .io_en_1( io_VwirePorts_3_17_4_en ),
       .io_en_0( io_VwirePorts_2_17_4_en ),
       .io_out( Vwire_63_io_out )
  );
  Vwire_0 Vwire_64(
       .io_in_1( io_VwirePorts_3_18_4_in ),
       .io_in_0( io_VwirePorts_2_18_4_in ),
       .io_en_1( io_VwirePorts_3_18_4_en ),
       .io_en_0( io_VwirePorts_2_18_4_en ),
       .io_out( Vwire_64_io_out )
  );
  Vwire_0 Vwire_65(
       .io_in_1( io_VwirePorts_3_19_4_in ),
       .io_in_0( io_VwirePorts_2_19_4_in ),
       .io_en_1( io_VwirePorts_3_19_4_en ),
       .io_en_0( io_VwirePorts_2_19_4_en ),
       .io_out( Vwire_65_io_out )
  );
  Vwire_0 Vwire_66(
       .io_in_1( io_VwirePorts_3_20_4_in ),
       .io_in_0( io_VwirePorts_2_20_4_in ),
       .io_en_1( io_VwirePorts_3_20_4_en ),
       .io_en_0( io_VwirePorts_2_20_4_en ),
       .io_out( Vwire_66_io_out )
  );
  Vwire_0 Vwire_67(
       .io_in_1( io_VwirePorts_3_21_4_in ),
       .io_in_0( io_VwirePorts_2_21_4_in ),
       .io_en_1( io_VwirePorts_3_21_4_en ),
       .io_en_0( io_VwirePorts_2_21_4_en ),
       .io_out( Vwire_67_io_out )
  );
  Vwire_0 Vwire_68(
       .io_in_1( io_VwirePorts_3_22_4_in ),
       .io_in_0( io_VwirePorts_2_22_4_in ),
       .io_en_1( io_VwirePorts_3_22_4_en ),
       .io_en_0( io_VwirePorts_2_22_4_en ),
       .io_out( Vwire_68_io_out )
  );
  Vwire_0 Vwire_69(
       .io_in_1( io_VwirePorts_1_0_4_in ),
       .io_in_0( io_VwirePorts_0_0_4_in ),
       .io_en_1( io_VwirePorts_1_0_4_en ),
       .io_en_0( io_VwirePorts_0_0_4_en ),
       .io_out( Vwire_69_io_out )
  );
  Vwire_0 Vwire_70(
       .io_in_1( io_VwirePorts_1_1_4_in ),
       .io_in_0( io_VwirePorts_0_1_4_in ),
       .io_en_1( io_VwirePorts_1_1_4_en ),
       .io_en_0( io_VwirePorts_0_1_4_en ),
       .io_out( Vwire_70_io_out )
  );
  Vwire_0 Vwire_71(
       .io_in_1( io_VwirePorts_1_2_4_in ),
       .io_in_0( io_VwirePorts_0_2_4_in ),
       .io_en_1( io_VwirePorts_1_2_4_en ),
       .io_en_0( io_VwirePorts_0_2_4_en ),
       .io_out( Vwire_71_io_out )
  );
  Vwire_0 Vwire_72(
       .io_in_1( io_VwirePorts_1_3_4_in ),
       .io_in_0( io_VwirePorts_0_3_4_in ),
       .io_en_1( io_VwirePorts_1_3_4_en ),
       .io_en_0( io_VwirePorts_0_3_4_en ),
       .io_out( Vwire_72_io_out )
  );
  Vwire_0 Vwire_73(
       .io_in_1( io_VwirePorts_1_4_4_in ),
       .io_in_0( io_VwirePorts_0_4_4_in ),
       .io_en_1( io_VwirePorts_1_4_4_en ),
       .io_en_0( io_VwirePorts_0_4_4_en ),
       .io_out( Vwire_73_io_out )
  );
  Vwire_0 Vwire_74(
       .io_in_1( io_VwirePorts_1_5_4_in ),
       .io_in_0( io_VwirePorts_0_5_4_in ),
       .io_en_1( io_VwirePorts_1_5_4_en ),
       .io_en_0( io_VwirePorts_0_5_4_en ),
       .io_out( Vwire_74_io_out )
  );
  Vwire_0 Vwire_75(
       .io_in_1( io_VwirePorts_1_6_4_in ),
       .io_in_0( io_VwirePorts_0_6_4_in ),
       .io_en_1( io_VwirePorts_1_6_4_en ),
       .io_en_0( io_VwirePorts_0_6_4_en ),
       .io_out( Vwire_75_io_out )
  );
  Vwire_0 Vwire_76(
       .io_in_1( io_VwirePorts_1_7_4_in ),
       .io_in_0( io_VwirePorts_0_7_4_in ),
       .io_en_1( io_VwirePorts_1_7_4_en ),
       .io_en_0( io_VwirePorts_0_7_4_en ),
       .io_out( Vwire_76_io_out )
  );
  Vwire_0 Vwire_77(
       .io_in_1( io_VwirePorts_1_8_4_in ),
       .io_in_0( io_VwirePorts_0_8_4_in ),
       .io_en_1( io_VwirePorts_1_8_4_en ),
       .io_en_0( io_VwirePorts_0_8_4_en ),
       .io_out( Vwire_77_io_out )
  );
  Vwire_0 Vwire_78(
       .io_in_1( io_VwirePorts_1_9_4_in ),
       .io_in_0( io_VwirePorts_0_9_4_in ),
       .io_en_1( io_VwirePorts_1_9_4_en ),
       .io_en_0( io_VwirePorts_0_9_4_en ),
       .io_out( Vwire_78_io_out )
  );
  Vwire_0 Vwire_79(
       .io_in_1( io_VwirePorts_1_10_4_in ),
       .io_in_0( io_VwirePorts_0_10_4_in ),
       .io_en_1( io_VwirePorts_1_10_4_en ),
       .io_en_0( io_VwirePorts_0_10_4_en ),
       .io_out( Vwire_79_io_out )
  );
  Vwire_0 Vwire_80(
       .io_in_1( io_VwirePorts_1_11_4_in ),
       .io_in_0( io_VwirePorts_0_11_4_in ),
       .io_en_1( io_VwirePorts_1_11_4_en ),
       .io_en_0( io_VwirePorts_0_11_4_en ),
       .io_out( Vwire_80_io_out )
  );
  Vwire_0 Vwire_81(
       .io_in_1( io_VwirePorts_1_12_4_in ),
       .io_in_0( io_VwirePorts_0_12_4_in ),
       .io_en_1( io_VwirePorts_1_12_4_en ),
       .io_en_0( io_VwirePorts_0_12_4_en ),
       .io_out( Vwire_81_io_out )
  );
  Vwire_0 Vwire_82(
       .io_in_1( io_VwirePorts_1_13_4_in ),
       .io_in_0( io_VwirePorts_0_13_4_in ),
       .io_en_1( io_VwirePorts_1_13_4_en ),
       .io_en_0( io_VwirePorts_0_13_4_en ),
       .io_out( Vwire_82_io_out )
  );
  Vwire_0 Vwire_83(
       .io_in_1( io_VwirePorts_1_14_4_in ),
       .io_in_0( io_VwirePorts_0_14_4_in ),
       .io_en_1( io_VwirePorts_1_14_4_en ),
       .io_en_0( io_VwirePorts_0_14_4_en ),
       .io_out( Vwire_83_io_out )
  );
  Vwire_0 Vwire_84(
       .io_in_1( io_VwirePorts_1_15_4_in ),
       .io_in_0( io_VwirePorts_0_15_4_in ),
       .io_en_1( io_VwirePorts_1_15_4_en ),
       .io_en_0( io_VwirePorts_0_15_4_en ),
       .io_out( Vwire_84_io_out )
  );
  Vwire_0 Vwire_85(
       .io_in_1( io_VwirePorts_1_16_4_in ),
       .io_in_0( io_VwirePorts_0_16_4_in ),
       .io_en_1( io_VwirePorts_1_16_4_en ),
       .io_en_0( io_VwirePorts_0_16_4_en ),
       .io_out( Vwire_85_io_out )
  );
  Vwire_0 Vwire_86(
       .io_in_1( io_VwirePorts_1_17_4_in ),
       .io_in_0( io_VwirePorts_0_17_4_in ),
       .io_en_1( io_VwirePorts_1_17_4_en ),
       .io_en_0( io_VwirePorts_0_17_4_en ),
       .io_out( Vwire_86_io_out )
  );
  Vwire_0 Vwire_87(
       .io_in_1( io_VwirePorts_1_18_4_in ),
       .io_in_0( io_VwirePorts_0_18_4_in ),
       .io_en_1( io_VwirePorts_1_18_4_en ),
       .io_en_0( io_VwirePorts_0_18_4_en ),
       .io_out( Vwire_87_io_out )
  );
  Vwire_0 Vwire_88(
       .io_in_1( io_VwirePorts_1_19_4_in ),
       .io_in_0( io_VwirePorts_0_19_4_in ),
       .io_en_1( io_VwirePorts_1_19_4_en ),
       .io_en_0( io_VwirePorts_0_19_4_en ),
       .io_out( Vwire_88_io_out )
  );
  Vwire_0 Vwire_89(
       .io_in_1( io_VwirePorts_1_20_4_in ),
       .io_in_0( io_VwirePorts_0_20_4_in ),
       .io_en_1( io_VwirePorts_1_20_4_en ),
       .io_en_0( io_VwirePorts_0_20_4_en ),
       .io_out( Vwire_89_io_out )
  );
  Vwire_0 Vwire_90(
       .io_in_1( io_VwirePorts_1_21_4_in ),
       .io_in_0( io_VwirePorts_0_21_4_in ),
       .io_en_1( io_VwirePorts_1_21_4_en ),
       .io_en_0( io_VwirePorts_0_21_4_en ),
       .io_out( Vwire_90_io_out )
  );
  Vwire_0 Vwire_91(
       .io_in_1( io_VwirePorts_1_22_4_in ),
       .io_in_0( io_VwirePorts_0_22_4_in ),
       .io_en_1( io_VwirePorts_1_22_4_en ),
       .io_en_0( io_VwirePorts_0_22_4_en ),
       .io_out( Vwire_91_io_out )
  );
  Vwire_1 Vwire_92(
       .io_in_2( io_VwirePorts_3_0_3_in ),
       .io_in_1( io_VwirePorts_2_0_3_in ),
       .io_in_0( io_VwirePorts_1_0_2_in ),
       .io_en_2( io_VwirePorts_3_0_3_en ),
       .io_en_1( io_VwirePorts_2_0_3_en ),
       .io_en_0( io_VwirePorts_1_0_2_en ),
       .io_out( Vwire_92_io_out )
  );
  Vwire_1 Vwire_93(
       .io_in_2( io_VwirePorts_3_1_3_in ),
       .io_in_1( io_VwirePorts_2_1_3_in ),
       .io_in_0( io_VwirePorts_1_1_2_in ),
       .io_en_2( io_VwirePorts_3_1_3_en ),
       .io_en_1( io_VwirePorts_2_1_3_en ),
       .io_en_0( io_VwirePorts_1_1_2_en ),
       .io_out( Vwire_93_io_out )
  );
  Vwire_1 Vwire_94(
       .io_in_2( io_VwirePorts_3_2_3_in ),
       .io_in_1( io_VwirePorts_2_2_3_in ),
       .io_in_0( io_VwirePorts_1_2_2_in ),
       .io_en_2( io_VwirePorts_3_2_3_en ),
       .io_en_1( io_VwirePorts_2_2_3_en ),
       .io_en_0( io_VwirePorts_1_2_2_en ),
       .io_out( Vwire_94_io_out )
  );
  Vwire_1 Vwire_95(
       .io_in_2( io_VwirePorts_3_3_3_in ),
       .io_in_1( io_VwirePorts_2_3_3_in ),
       .io_in_0( io_VwirePorts_1_3_2_in ),
       .io_en_2( io_VwirePorts_3_3_3_en ),
       .io_en_1( io_VwirePorts_2_3_3_en ),
       .io_en_0( io_VwirePorts_1_3_2_en ),
       .io_out( Vwire_95_io_out )
  );
  Vwire_1 Vwire_96(
       .io_in_2( io_VwirePorts_3_4_3_in ),
       .io_in_1( io_VwirePorts_2_4_3_in ),
       .io_in_0( io_VwirePorts_1_4_2_in ),
       .io_en_2( io_VwirePorts_3_4_3_en ),
       .io_en_1( io_VwirePorts_2_4_3_en ),
       .io_en_0( io_VwirePorts_1_4_2_en ),
       .io_out( Vwire_96_io_out )
  );
  Vwire_1 Vwire_97(
       .io_in_2( io_VwirePorts_3_5_3_in ),
       .io_in_1( io_VwirePorts_2_5_3_in ),
       .io_in_0( io_VwirePorts_1_5_2_in ),
       .io_en_2( io_VwirePorts_3_5_3_en ),
       .io_en_1( io_VwirePorts_2_5_3_en ),
       .io_en_0( io_VwirePorts_1_5_2_en ),
       .io_out( Vwire_97_io_out )
  );
  Vwire_1 Vwire_98(
       .io_in_2( io_VwirePorts_3_6_3_in ),
       .io_in_1( io_VwirePorts_2_6_3_in ),
       .io_in_0( io_VwirePorts_1_6_2_in ),
       .io_en_2( io_VwirePorts_3_6_3_en ),
       .io_en_1( io_VwirePorts_2_6_3_en ),
       .io_en_0( io_VwirePorts_1_6_2_en ),
       .io_out( Vwire_98_io_out )
  );
  Vwire_1 Vwire_99(
       .io_in_2( io_VwirePorts_3_7_3_in ),
       .io_in_1( io_VwirePorts_2_7_3_in ),
       .io_in_0( io_VwirePorts_1_7_2_in ),
       .io_en_2( io_VwirePorts_3_7_3_en ),
       .io_en_1( io_VwirePorts_2_7_3_en ),
       .io_en_0( io_VwirePorts_1_7_2_en ),
       .io_out( Vwire_99_io_out )
  );
  Vwire_1 Vwire_100(
       .io_in_2( io_VwirePorts_3_8_3_in ),
       .io_in_1( io_VwirePorts_2_8_3_in ),
       .io_in_0( io_VwirePorts_1_8_2_in ),
       .io_en_2( io_VwirePorts_3_8_3_en ),
       .io_en_1( io_VwirePorts_2_8_3_en ),
       .io_en_0( io_VwirePorts_1_8_2_en ),
       .io_out( Vwire_100_io_out )
  );
  Vwire_1 Vwire_101(
       .io_in_2( io_VwirePorts_3_9_3_in ),
       .io_in_1( io_VwirePorts_2_9_3_in ),
       .io_in_0( io_VwirePorts_1_9_2_in ),
       .io_en_2( io_VwirePorts_3_9_3_en ),
       .io_en_1( io_VwirePorts_2_9_3_en ),
       .io_en_0( io_VwirePorts_1_9_2_en ),
       .io_out( Vwire_101_io_out )
  );
  Vwire_1 Vwire_102(
       .io_in_2( io_VwirePorts_3_10_3_in ),
       .io_in_1( io_VwirePorts_2_10_3_in ),
       .io_in_0( io_VwirePorts_1_10_2_in ),
       .io_en_2( io_VwirePorts_3_10_3_en ),
       .io_en_1( io_VwirePorts_2_10_3_en ),
       .io_en_0( io_VwirePorts_1_10_2_en ),
       .io_out( Vwire_102_io_out )
  );
  Vwire_1 Vwire_103(
       .io_in_2( io_VwirePorts_3_11_3_in ),
       .io_in_1( io_VwirePorts_2_11_3_in ),
       .io_in_0( io_VwirePorts_1_11_2_in ),
       .io_en_2( io_VwirePorts_3_11_3_en ),
       .io_en_1( io_VwirePorts_2_11_3_en ),
       .io_en_0( io_VwirePorts_1_11_2_en ),
       .io_out( Vwire_103_io_out )
  );
  Vwire_1 Vwire_104(
       .io_in_2( io_VwirePorts_3_12_3_in ),
       .io_in_1( io_VwirePorts_2_12_3_in ),
       .io_in_0( io_VwirePorts_1_12_2_in ),
       .io_en_2( io_VwirePorts_3_12_3_en ),
       .io_en_1( io_VwirePorts_2_12_3_en ),
       .io_en_0( io_VwirePorts_1_12_2_en ),
       .io_out( Vwire_104_io_out )
  );
  Vwire_1 Vwire_105(
       .io_in_2( io_VwirePorts_3_13_3_in ),
       .io_in_1( io_VwirePorts_2_13_3_in ),
       .io_in_0( io_VwirePorts_1_13_2_in ),
       .io_en_2( io_VwirePorts_3_13_3_en ),
       .io_en_1( io_VwirePorts_2_13_3_en ),
       .io_en_0( io_VwirePorts_1_13_2_en ),
       .io_out( Vwire_105_io_out )
  );
  Vwire_1 Vwire_106(
       .io_in_2( io_VwirePorts_3_14_3_in ),
       .io_in_1( io_VwirePorts_2_14_3_in ),
       .io_in_0( io_VwirePorts_1_14_2_in ),
       .io_en_2( io_VwirePorts_3_14_3_en ),
       .io_en_1( io_VwirePorts_2_14_3_en ),
       .io_en_0( io_VwirePorts_1_14_2_en ),
       .io_out( Vwire_106_io_out )
  );
  Vwire_1 Vwire_107(
       .io_in_2( io_VwirePorts_3_15_3_in ),
       .io_in_1( io_VwirePorts_2_15_3_in ),
       .io_in_0( io_VwirePorts_1_15_2_in ),
       .io_en_2( io_VwirePorts_3_15_3_en ),
       .io_en_1( io_VwirePorts_2_15_3_en ),
       .io_en_0( io_VwirePorts_1_15_2_en ),
       .io_out( Vwire_107_io_out )
  );
  Vwire_1 Vwire_108(
       .io_in_2( io_VwirePorts_3_16_3_in ),
       .io_in_1( io_VwirePorts_2_16_3_in ),
       .io_in_0( io_VwirePorts_1_16_2_in ),
       .io_en_2( io_VwirePorts_3_16_3_en ),
       .io_en_1( io_VwirePorts_2_16_3_en ),
       .io_en_0( io_VwirePorts_1_16_2_en ),
       .io_out( Vwire_108_io_out )
  );
  Vwire_1 Vwire_109(
       .io_in_2( io_VwirePorts_3_17_3_in ),
       .io_in_1( io_VwirePorts_2_17_3_in ),
       .io_in_0( io_VwirePorts_1_17_2_in ),
       .io_en_2( io_VwirePorts_3_17_3_en ),
       .io_en_1( io_VwirePorts_2_17_3_en ),
       .io_en_0( io_VwirePorts_1_17_2_en ),
       .io_out( Vwire_109_io_out )
  );
  Vwire_1 Vwire_110(
       .io_in_2( io_VwirePorts_3_18_3_in ),
       .io_in_1( io_VwirePorts_2_18_3_in ),
       .io_in_0( io_VwirePorts_1_18_2_in ),
       .io_en_2( io_VwirePorts_3_18_3_en ),
       .io_en_1( io_VwirePorts_2_18_3_en ),
       .io_en_0( io_VwirePorts_1_18_2_en ),
       .io_out( Vwire_110_io_out )
  );
  Vwire_1 Vwire_111(
       .io_in_2( io_VwirePorts_3_19_3_in ),
       .io_in_1( io_VwirePorts_2_19_3_in ),
       .io_in_0( io_VwirePorts_1_19_2_in ),
       .io_en_2( io_VwirePorts_3_19_3_en ),
       .io_en_1( io_VwirePorts_2_19_3_en ),
       .io_en_0( io_VwirePorts_1_19_2_en ),
       .io_out( Vwire_111_io_out )
  );
  Vwire_1 Vwire_112(
       .io_in_2( io_VwirePorts_3_20_3_in ),
       .io_in_1( io_VwirePorts_2_20_3_in ),
       .io_in_0( io_VwirePorts_1_20_2_in ),
       .io_en_2( io_VwirePorts_3_20_3_en ),
       .io_en_1( io_VwirePorts_2_20_3_en ),
       .io_en_0( io_VwirePorts_1_20_2_en ),
       .io_out( Vwire_112_io_out )
  );
  Vwire_1 Vwire_113(
       .io_in_2( io_VwirePorts_3_21_3_in ),
       .io_in_1( io_VwirePorts_2_21_3_in ),
       .io_in_0( io_VwirePorts_1_21_2_in ),
       .io_en_2( io_VwirePorts_3_21_3_en ),
       .io_en_1( io_VwirePorts_2_21_3_en ),
       .io_en_0( io_VwirePorts_1_21_2_en ),
       .io_out( Vwire_113_io_out )
  );
  Vwire_1 Vwire_114(
       .io_in_2( io_VwirePorts_3_22_3_in ),
       .io_in_1( io_VwirePorts_2_22_3_in ),
       .io_in_0( io_VwirePorts_1_22_2_in ),
       .io_en_2( io_VwirePorts_3_22_3_en ),
       .io_en_1( io_VwirePorts_2_22_3_en ),
       .io_en_0( io_VwirePorts_1_22_2_en ),
       .io_out( Vwire_114_io_out )
  );
  Vwire_1 Vwire_115(
       .io_in_2( io_VwirePorts_2_0_2_in ),
       .io_in_1( io_VwirePorts_1_0_3_in ),
       .io_in_0( io_VwirePorts_0_0_3_in ),
       .io_en_2( io_VwirePorts_2_0_2_en ),
       .io_en_1( io_VwirePorts_1_0_3_en ),
       .io_en_0( io_VwirePorts_0_0_3_en ),
       .io_out( Vwire_115_io_out )
  );
  Vwire_1 Vwire_116(
       .io_in_2( io_VwirePorts_2_1_2_in ),
       .io_in_1( io_VwirePorts_1_1_3_in ),
       .io_in_0( io_VwirePorts_0_1_3_in ),
       .io_en_2( io_VwirePorts_2_1_2_en ),
       .io_en_1( io_VwirePorts_1_1_3_en ),
       .io_en_0( io_VwirePorts_0_1_3_en ),
       .io_out( Vwire_116_io_out )
  );
  Vwire_1 Vwire_117(
       .io_in_2( io_VwirePorts_2_2_2_in ),
       .io_in_1( io_VwirePorts_1_2_3_in ),
       .io_in_0( io_VwirePorts_0_2_3_in ),
       .io_en_2( io_VwirePorts_2_2_2_en ),
       .io_en_1( io_VwirePorts_1_2_3_en ),
       .io_en_0( io_VwirePorts_0_2_3_en ),
       .io_out( Vwire_117_io_out )
  );
  Vwire_1 Vwire_118(
       .io_in_2( io_VwirePorts_2_3_2_in ),
       .io_in_1( io_VwirePorts_1_3_3_in ),
       .io_in_0( io_VwirePorts_0_3_3_in ),
       .io_en_2( io_VwirePorts_2_3_2_en ),
       .io_en_1( io_VwirePorts_1_3_3_en ),
       .io_en_0( io_VwirePorts_0_3_3_en ),
       .io_out( Vwire_118_io_out )
  );
  Vwire_1 Vwire_119(
       .io_in_2( io_VwirePorts_2_4_2_in ),
       .io_in_1( io_VwirePorts_1_4_3_in ),
       .io_in_0( io_VwirePorts_0_4_3_in ),
       .io_en_2( io_VwirePorts_2_4_2_en ),
       .io_en_1( io_VwirePorts_1_4_3_en ),
       .io_en_0( io_VwirePorts_0_4_3_en ),
       .io_out( Vwire_119_io_out )
  );
  Vwire_1 Vwire_120(
       .io_in_2( io_VwirePorts_2_5_2_in ),
       .io_in_1( io_VwirePorts_1_5_3_in ),
       .io_in_0( io_VwirePorts_0_5_3_in ),
       .io_en_2( io_VwirePorts_2_5_2_en ),
       .io_en_1( io_VwirePorts_1_5_3_en ),
       .io_en_0( io_VwirePorts_0_5_3_en ),
       .io_out( Vwire_120_io_out )
  );
  Vwire_1 Vwire_121(
       .io_in_2( io_VwirePorts_2_6_2_in ),
       .io_in_1( io_VwirePorts_1_6_3_in ),
       .io_in_0( io_VwirePorts_0_6_3_in ),
       .io_en_2( io_VwirePorts_2_6_2_en ),
       .io_en_1( io_VwirePorts_1_6_3_en ),
       .io_en_0( io_VwirePorts_0_6_3_en ),
       .io_out( Vwire_121_io_out )
  );
  Vwire_1 Vwire_122(
       .io_in_2( io_VwirePorts_2_7_2_in ),
       .io_in_1( io_VwirePorts_1_7_3_in ),
       .io_in_0( io_VwirePorts_0_7_3_in ),
       .io_en_2( io_VwirePorts_2_7_2_en ),
       .io_en_1( io_VwirePorts_1_7_3_en ),
       .io_en_0( io_VwirePorts_0_7_3_en ),
       .io_out( Vwire_122_io_out )
  );
  Vwire_1 Vwire_123(
       .io_in_2( io_VwirePorts_2_8_2_in ),
       .io_in_1( io_VwirePorts_1_8_3_in ),
       .io_in_0( io_VwirePorts_0_8_3_in ),
       .io_en_2( io_VwirePorts_2_8_2_en ),
       .io_en_1( io_VwirePorts_1_8_3_en ),
       .io_en_0( io_VwirePorts_0_8_3_en ),
       .io_out( Vwire_123_io_out )
  );
  Vwire_1 Vwire_124(
       .io_in_2( io_VwirePorts_2_9_2_in ),
       .io_in_1( io_VwirePorts_1_9_3_in ),
       .io_in_0( io_VwirePorts_0_9_3_in ),
       .io_en_2( io_VwirePorts_2_9_2_en ),
       .io_en_1( io_VwirePorts_1_9_3_en ),
       .io_en_0( io_VwirePorts_0_9_3_en ),
       .io_out( Vwire_124_io_out )
  );
  Vwire_1 Vwire_125(
       .io_in_2( io_VwirePorts_2_10_2_in ),
       .io_in_1( io_VwirePorts_1_10_3_in ),
       .io_in_0( io_VwirePorts_0_10_3_in ),
       .io_en_2( io_VwirePorts_2_10_2_en ),
       .io_en_1( io_VwirePorts_1_10_3_en ),
       .io_en_0( io_VwirePorts_0_10_3_en ),
       .io_out( Vwire_125_io_out )
  );
  Vwire_1 Vwire_126(
       .io_in_2( io_VwirePorts_2_11_2_in ),
       .io_in_1( io_VwirePorts_1_11_3_in ),
       .io_in_0( io_VwirePorts_0_11_3_in ),
       .io_en_2( io_VwirePorts_2_11_2_en ),
       .io_en_1( io_VwirePorts_1_11_3_en ),
       .io_en_0( io_VwirePorts_0_11_3_en ),
       .io_out( Vwire_126_io_out )
  );
  Vwire_1 Vwire_127(
       .io_in_2( io_VwirePorts_2_12_2_in ),
       .io_in_1( io_VwirePorts_1_12_3_in ),
       .io_in_0( io_VwirePorts_0_12_3_in ),
       .io_en_2( io_VwirePorts_2_12_2_en ),
       .io_en_1( io_VwirePorts_1_12_3_en ),
       .io_en_0( io_VwirePorts_0_12_3_en ),
       .io_out( Vwire_127_io_out )
  );
  Vwire_1 Vwire_128(
       .io_in_2( io_VwirePorts_2_13_2_in ),
       .io_in_1( io_VwirePorts_1_13_3_in ),
       .io_in_0( io_VwirePorts_0_13_3_in ),
       .io_en_2( io_VwirePorts_2_13_2_en ),
       .io_en_1( io_VwirePorts_1_13_3_en ),
       .io_en_0( io_VwirePorts_0_13_3_en ),
       .io_out( Vwire_128_io_out )
  );
  Vwire_1 Vwire_129(
       .io_in_2( io_VwirePorts_2_14_2_in ),
       .io_in_1( io_VwirePorts_1_14_3_in ),
       .io_in_0( io_VwirePorts_0_14_3_in ),
       .io_en_2( io_VwirePorts_2_14_2_en ),
       .io_en_1( io_VwirePorts_1_14_3_en ),
       .io_en_0( io_VwirePorts_0_14_3_en ),
       .io_out( Vwire_129_io_out )
  );
  Vwire_1 Vwire_130(
       .io_in_2( io_VwirePorts_2_15_2_in ),
       .io_in_1( io_VwirePorts_1_15_3_in ),
       .io_in_0( io_VwirePorts_0_15_3_in ),
       .io_en_2( io_VwirePorts_2_15_2_en ),
       .io_en_1( io_VwirePorts_1_15_3_en ),
       .io_en_0( io_VwirePorts_0_15_3_en ),
       .io_out( Vwire_130_io_out )
  );
  Vwire_1 Vwire_131(
       .io_in_2( io_VwirePorts_2_16_2_in ),
       .io_in_1( io_VwirePorts_1_16_3_in ),
       .io_in_0( io_VwirePorts_0_16_3_in ),
       .io_en_2( io_VwirePorts_2_16_2_en ),
       .io_en_1( io_VwirePorts_1_16_3_en ),
       .io_en_0( io_VwirePorts_0_16_3_en ),
       .io_out( Vwire_131_io_out )
  );
  Vwire_1 Vwire_132(
       .io_in_2( io_VwirePorts_2_17_2_in ),
       .io_in_1( io_VwirePorts_1_17_3_in ),
       .io_in_0( io_VwirePorts_0_17_3_in ),
       .io_en_2( io_VwirePorts_2_17_2_en ),
       .io_en_1( io_VwirePorts_1_17_3_en ),
       .io_en_0( io_VwirePorts_0_17_3_en ),
       .io_out( Vwire_132_io_out )
  );
  Vwire_1 Vwire_133(
       .io_in_2( io_VwirePorts_2_18_2_in ),
       .io_in_1( io_VwirePorts_1_18_3_in ),
       .io_in_0( io_VwirePorts_0_18_3_in ),
       .io_en_2( io_VwirePorts_2_18_2_en ),
       .io_en_1( io_VwirePorts_1_18_3_en ),
       .io_en_0( io_VwirePorts_0_18_3_en ),
       .io_out( Vwire_133_io_out )
  );
  Vwire_1 Vwire_134(
       .io_in_2( io_VwirePorts_2_19_2_in ),
       .io_in_1( io_VwirePorts_1_19_3_in ),
       .io_in_0( io_VwirePorts_0_19_3_in ),
       .io_en_2( io_VwirePorts_2_19_2_en ),
       .io_en_1( io_VwirePorts_1_19_3_en ),
       .io_en_0( io_VwirePorts_0_19_3_en ),
       .io_out( Vwire_134_io_out )
  );
  Vwire_1 Vwire_135(
       .io_in_2( io_VwirePorts_2_20_2_in ),
       .io_in_1( io_VwirePorts_1_20_3_in ),
       .io_in_0( io_VwirePorts_0_20_3_in ),
       .io_en_2( io_VwirePorts_2_20_2_en ),
       .io_en_1( io_VwirePorts_1_20_3_en ),
       .io_en_0( io_VwirePorts_0_20_3_en ),
       .io_out( Vwire_135_io_out )
  );
  Vwire_1 Vwire_136(
       .io_in_2( io_VwirePorts_2_21_2_in ),
       .io_in_1( io_VwirePorts_1_21_3_in ),
       .io_in_0( io_VwirePorts_0_21_3_in ),
       .io_en_2( io_VwirePorts_2_21_2_en ),
       .io_en_1( io_VwirePorts_1_21_3_en ),
       .io_en_0( io_VwirePorts_0_21_3_en ),
       .io_out( Vwire_136_io_out )
  );
  Vwire_1 Vwire_137(
       .io_in_2( io_VwirePorts_2_22_2_in ),
       .io_in_1( io_VwirePorts_1_22_3_in ),
       .io_in_0( io_VwirePorts_0_22_3_in ),
       .io_en_2( io_VwirePorts_2_22_2_en ),
       .io_en_1( io_VwirePorts_1_22_3_en ),
       .io_en_0( io_VwirePorts_0_22_3_en ),
       .io_out( Vwire_137_io_out )
  );
  Vwire_2 Vwire_138(
       .io_in_3( io_VwirePorts_3_0_0_in ),
       .io_in_2( io_VwirePorts_2_0_1_in ),
       .io_in_1( io_VwirePorts_1_0_1_in ),
       .io_in_0( io_VwirePorts_0_0_0_in ),
       .io_en_3( io_VwirePorts_3_0_0_en ),
       .io_en_2( io_VwirePorts_2_0_1_en ),
       .io_en_1( io_VwirePorts_1_0_1_en ),
       .io_en_0( io_VwirePorts_0_0_0_en ),
       .io_out( Vwire_138_io_out )
  );
  Vwire_2 Vwire_139(
       .io_in_3( io_VwirePorts_3_1_0_in ),
       .io_in_2( io_VwirePorts_2_1_1_in ),
       .io_in_1( io_VwirePorts_1_1_1_in ),
       .io_in_0( io_VwirePorts_0_1_0_in ),
       .io_en_3( io_VwirePorts_3_1_0_en ),
       .io_en_2( io_VwirePorts_2_1_1_en ),
       .io_en_1( io_VwirePorts_1_1_1_en ),
       .io_en_0( io_VwirePorts_0_1_0_en ),
       .io_out( Vwire_139_io_out )
  );
  Vwire_2 Vwire_140(
       .io_in_3( io_VwirePorts_3_2_0_in ),
       .io_in_2( io_VwirePorts_2_2_1_in ),
       .io_in_1( io_VwirePorts_1_2_1_in ),
       .io_in_0( io_VwirePorts_0_2_0_in ),
       .io_en_3( io_VwirePorts_3_2_0_en ),
       .io_en_2( io_VwirePorts_2_2_1_en ),
       .io_en_1( io_VwirePorts_1_2_1_en ),
       .io_en_0( io_VwirePorts_0_2_0_en ),
       .io_out( Vwire_140_io_out )
  );
  Vwire_2 Vwire_141(
       .io_in_3( io_VwirePorts_3_3_0_in ),
       .io_in_2( io_VwirePorts_2_3_1_in ),
       .io_in_1( io_VwirePorts_1_3_1_in ),
       .io_in_0( io_VwirePorts_0_3_0_in ),
       .io_en_3( io_VwirePorts_3_3_0_en ),
       .io_en_2( io_VwirePorts_2_3_1_en ),
       .io_en_1( io_VwirePorts_1_3_1_en ),
       .io_en_0( io_VwirePorts_0_3_0_en ),
       .io_out( Vwire_141_io_out )
  );
  Vwire_2 Vwire_142(
       .io_in_3( io_VwirePorts_3_4_0_in ),
       .io_in_2( io_VwirePorts_2_4_1_in ),
       .io_in_1( io_VwirePorts_1_4_1_in ),
       .io_in_0( io_VwirePorts_0_4_0_in ),
       .io_en_3( io_VwirePorts_3_4_0_en ),
       .io_en_2( io_VwirePorts_2_4_1_en ),
       .io_en_1( io_VwirePorts_1_4_1_en ),
       .io_en_0( io_VwirePorts_0_4_0_en ),
       .io_out( Vwire_142_io_out )
  );
  Vwire_2 Vwire_143(
       .io_in_3( io_VwirePorts_3_5_0_in ),
       .io_in_2( io_VwirePorts_2_5_1_in ),
       .io_in_1( io_VwirePorts_1_5_1_in ),
       .io_in_0( io_VwirePorts_0_5_0_in ),
       .io_en_3( io_VwirePorts_3_5_0_en ),
       .io_en_2( io_VwirePorts_2_5_1_en ),
       .io_en_1( io_VwirePorts_1_5_1_en ),
       .io_en_0( io_VwirePorts_0_5_0_en ),
       .io_out( Vwire_143_io_out )
  );
  Vwire_2 Vwire_144(
       .io_in_3( io_VwirePorts_3_6_0_in ),
       .io_in_2( io_VwirePorts_2_6_1_in ),
       .io_in_1( io_VwirePorts_1_6_1_in ),
       .io_in_0( io_VwirePorts_0_6_0_in ),
       .io_en_3( io_VwirePorts_3_6_0_en ),
       .io_en_2( io_VwirePorts_2_6_1_en ),
       .io_en_1( io_VwirePorts_1_6_1_en ),
       .io_en_0( io_VwirePorts_0_6_0_en ),
       .io_out( Vwire_144_io_out )
  );
  Vwire_2 Vwire_145(
       .io_in_3( io_VwirePorts_3_7_0_in ),
       .io_in_2( io_VwirePorts_2_7_1_in ),
       .io_in_1( io_VwirePorts_1_7_1_in ),
       .io_in_0( io_VwirePorts_0_7_0_in ),
       .io_en_3( io_VwirePorts_3_7_0_en ),
       .io_en_2( io_VwirePorts_2_7_1_en ),
       .io_en_1( io_VwirePorts_1_7_1_en ),
       .io_en_0( io_VwirePorts_0_7_0_en ),
       .io_out( Vwire_145_io_out )
  );
  Vwire_2 Vwire_146(
       .io_in_3( io_VwirePorts_3_8_0_in ),
       .io_in_2( io_VwirePorts_2_8_1_in ),
       .io_in_1( io_VwirePorts_1_8_1_in ),
       .io_in_0( io_VwirePorts_0_8_0_in ),
       .io_en_3( io_VwirePorts_3_8_0_en ),
       .io_en_2( io_VwirePorts_2_8_1_en ),
       .io_en_1( io_VwirePorts_1_8_1_en ),
       .io_en_0( io_VwirePorts_0_8_0_en ),
       .io_out( Vwire_146_io_out )
  );
  Vwire_2 Vwire_147(
       .io_in_3( io_VwirePorts_3_9_0_in ),
       .io_in_2( io_VwirePorts_2_9_1_in ),
       .io_in_1( io_VwirePorts_1_9_1_in ),
       .io_in_0( io_VwirePorts_0_9_0_in ),
       .io_en_3( io_VwirePorts_3_9_0_en ),
       .io_en_2( io_VwirePorts_2_9_1_en ),
       .io_en_1( io_VwirePorts_1_9_1_en ),
       .io_en_0( io_VwirePorts_0_9_0_en ),
       .io_out( Vwire_147_io_out )
  );
  Vwire_2 Vwire_148(
       .io_in_3( io_VwirePorts_3_10_0_in ),
       .io_in_2( io_VwirePorts_2_10_1_in ),
       .io_in_1( io_VwirePorts_1_10_1_in ),
       .io_in_0( io_VwirePorts_0_10_0_in ),
       .io_en_3( io_VwirePorts_3_10_0_en ),
       .io_en_2( io_VwirePorts_2_10_1_en ),
       .io_en_1( io_VwirePorts_1_10_1_en ),
       .io_en_0( io_VwirePorts_0_10_0_en ),
       .io_out( Vwire_148_io_out )
  );
  Vwire_2 Vwire_149(
       .io_in_3( io_VwirePorts_3_11_0_in ),
       .io_in_2( io_VwirePorts_2_11_1_in ),
       .io_in_1( io_VwirePorts_1_11_1_in ),
       .io_in_0( io_VwirePorts_0_11_0_in ),
       .io_en_3( io_VwirePorts_3_11_0_en ),
       .io_en_2( io_VwirePorts_2_11_1_en ),
       .io_en_1( io_VwirePorts_1_11_1_en ),
       .io_en_0( io_VwirePorts_0_11_0_en ),
       .io_out( Vwire_149_io_out )
  );
  Vwire_2 Vwire_150(
       .io_in_3( io_VwirePorts_3_12_0_in ),
       .io_in_2( io_VwirePorts_2_12_1_in ),
       .io_in_1( io_VwirePorts_1_12_1_in ),
       .io_in_0( io_VwirePorts_0_12_0_in ),
       .io_en_3( io_VwirePorts_3_12_0_en ),
       .io_en_2( io_VwirePorts_2_12_1_en ),
       .io_en_1( io_VwirePorts_1_12_1_en ),
       .io_en_0( io_VwirePorts_0_12_0_en ),
       .io_out( Vwire_150_io_out )
  );
  Vwire_2 Vwire_151(
       .io_in_3( io_VwirePorts_3_13_0_in ),
       .io_in_2( io_VwirePorts_2_13_1_in ),
       .io_in_1( io_VwirePorts_1_13_1_in ),
       .io_in_0( io_VwirePorts_0_13_0_in ),
       .io_en_3( io_VwirePorts_3_13_0_en ),
       .io_en_2( io_VwirePorts_2_13_1_en ),
       .io_en_1( io_VwirePorts_1_13_1_en ),
       .io_en_0( io_VwirePorts_0_13_0_en ),
       .io_out( Vwire_151_io_out )
  );
  Vwire_2 Vwire_152(
       .io_in_3( io_VwirePorts_3_14_0_in ),
       .io_in_2( io_VwirePorts_2_14_1_in ),
       .io_in_1( io_VwirePorts_1_14_1_in ),
       .io_in_0( io_VwirePorts_0_14_0_in ),
       .io_en_3( io_VwirePorts_3_14_0_en ),
       .io_en_2( io_VwirePorts_2_14_1_en ),
       .io_en_1( io_VwirePorts_1_14_1_en ),
       .io_en_0( io_VwirePorts_0_14_0_en ),
       .io_out( Vwire_152_io_out )
  );
  Vwire_2 Vwire_153(
       .io_in_3( io_VwirePorts_3_15_0_in ),
       .io_in_2( io_VwirePorts_2_15_1_in ),
       .io_in_1( io_VwirePorts_1_15_1_in ),
       .io_in_0( io_VwirePorts_0_15_0_in ),
       .io_en_3( io_VwirePorts_3_15_0_en ),
       .io_en_2( io_VwirePorts_2_15_1_en ),
       .io_en_1( io_VwirePorts_1_15_1_en ),
       .io_en_0( io_VwirePorts_0_15_0_en ),
       .io_out( Vwire_153_io_out )
  );
  Vwire_2 Vwire_154(
       .io_in_3( io_VwirePorts_3_16_0_in ),
       .io_in_2( io_VwirePorts_2_16_1_in ),
       .io_in_1( io_VwirePorts_1_16_1_in ),
       .io_in_0( io_VwirePorts_0_16_0_in ),
       .io_en_3( io_VwirePorts_3_16_0_en ),
       .io_en_2( io_VwirePorts_2_16_1_en ),
       .io_en_1( io_VwirePorts_1_16_1_en ),
       .io_en_0( io_VwirePorts_0_16_0_en ),
       .io_out( Vwire_154_io_out )
  );
  Vwire_2 Vwire_155(
       .io_in_3( io_VwirePorts_3_17_0_in ),
       .io_in_2( io_VwirePorts_2_17_1_in ),
       .io_in_1( io_VwirePorts_1_17_1_in ),
       .io_in_0( io_VwirePorts_0_17_0_in ),
       .io_en_3( io_VwirePorts_3_17_0_en ),
       .io_en_2( io_VwirePorts_2_17_1_en ),
       .io_en_1( io_VwirePorts_1_17_1_en ),
       .io_en_0( io_VwirePorts_0_17_0_en ),
       .io_out( Vwire_155_io_out )
  );
  Vwire_2 Vwire_156(
       .io_in_3( io_VwirePorts_3_18_0_in ),
       .io_in_2( io_VwirePorts_2_18_1_in ),
       .io_in_1( io_VwirePorts_1_18_1_in ),
       .io_in_0( io_VwirePorts_0_18_0_in ),
       .io_en_3( io_VwirePorts_3_18_0_en ),
       .io_en_2( io_VwirePorts_2_18_1_en ),
       .io_en_1( io_VwirePorts_1_18_1_en ),
       .io_en_0( io_VwirePorts_0_18_0_en ),
       .io_out( Vwire_156_io_out )
  );
  Vwire_2 Vwire_157(
       .io_in_3( io_VwirePorts_3_19_0_in ),
       .io_in_2( io_VwirePorts_2_19_1_in ),
       .io_in_1( io_VwirePorts_1_19_1_in ),
       .io_in_0( io_VwirePorts_0_19_0_in ),
       .io_en_3( io_VwirePorts_3_19_0_en ),
       .io_en_2( io_VwirePorts_2_19_1_en ),
       .io_en_1( io_VwirePorts_1_19_1_en ),
       .io_en_0( io_VwirePorts_0_19_0_en ),
       .io_out( Vwire_157_io_out )
  );
  Vwire_2 Vwire_158(
       .io_in_3( io_VwirePorts_3_20_0_in ),
       .io_in_2( io_VwirePorts_2_20_1_in ),
       .io_in_1( io_VwirePorts_1_20_1_in ),
       .io_in_0( io_VwirePorts_0_20_0_in ),
       .io_en_3( io_VwirePorts_3_20_0_en ),
       .io_en_2( io_VwirePorts_2_20_1_en ),
       .io_en_1( io_VwirePorts_1_20_1_en ),
       .io_en_0( io_VwirePorts_0_20_0_en ),
       .io_out( Vwire_158_io_out )
  );
  Vwire_2 Vwire_159(
       .io_in_3( io_VwirePorts_3_21_0_in ),
       .io_in_2( io_VwirePorts_2_21_1_in ),
       .io_in_1( io_VwirePorts_1_21_1_in ),
       .io_in_0( io_VwirePorts_0_21_0_in ),
       .io_en_3( io_VwirePorts_3_21_0_en ),
       .io_en_2( io_VwirePorts_2_21_1_en ),
       .io_en_1( io_VwirePorts_1_21_1_en ),
       .io_en_0( io_VwirePorts_0_21_0_en ),
       .io_out( Vwire_159_io_out )
  );
  Vwire_2 Vwire_160(
       .io_in_3( io_VwirePorts_3_22_0_in ),
       .io_in_2( io_VwirePorts_2_22_1_in ),
       .io_in_1( io_VwirePorts_1_22_1_in ),
       .io_in_0( io_VwirePorts_0_22_0_in ),
       .io_en_3( io_VwirePorts_3_22_0_en ),
       .io_en_2( io_VwirePorts_2_22_1_en ),
       .io_en_1( io_VwirePorts_1_22_1_en ),
       .io_en_0( io_VwirePorts_0_22_0_en ),
       .io_out( Vwire_160_io_out )
  );
  Vwire_2 Vwire_161(
       .io_in_3( io_VwirePorts_3_0_5_in ),
       .io_in_2( io_VwirePorts_2_0_5_in ),
       .io_in_1( io_VwirePorts_1_0_5_in ),
       .io_in_0( io_VwirePorts_0_0_5_in ),
       .io_en_3( io_VwirePorts_3_0_5_en ),
       .io_en_2( io_VwirePorts_2_0_5_en ),
       .io_en_1( io_VwirePorts_1_0_5_en ),
       .io_en_0( io_VwirePorts_0_0_5_en ),
       .io_out( Vwire_161_io_out )
  );
  Vwire_2 Vwire_162(
       .io_in_3( io_VwirePorts_3_1_5_in ),
       .io_in_2( io_VwirePorts_2_1_5_in ),
       .io_in_1( io_VwirePorts_1_1_5_in ),
       .io_in_0( io_VwirePorts_0_1_5_in ),
       .io_en_3( io_VwirePorts_3_1_5_en ),
       .io_en_2( io_VwirePorts_2_1_5_en ),
       .io_en_1( io_VwirePorts_1_1_5_en ),
       .io_en_0( io_VwirePorts_0_1_5_en ),
       .io_out( Vwire_162_io_out )
  );
  Vwire_2 Vwire_163(
       .io_in_3( io_VwirePorts_3_2_5_in ),
       .io_in_2( io_VwirePorts_2_2_5_in ),
       .io_in_1( io_VwirePorts_1_2_5_in ),
       .io_in_0( io_VwirePorts_0_2_5_in ),
       .io_en_3( io_VwirePorts_3_2_5_en ),
       .io_en_2( io_VwirePorts_2_2_5_en ),
       .io_en_1( io_VwirePorts_1_2_5_en ),
       .io_en_0( io_VwirePorts_0_2_5_en ),
       .io_out( Vwire_163_io_out )
  );
  Vwire_2 Vwire_164(
       .io_in_3( io_VwirePorts_3_3_5_in ),
       .io_in_2( io_VwirePorts_2_3_5_in ),
       .io_in_1( io_VwirePorts_1_3_5_in ),
       .io_in_0( io_VwirePorts_0_3_5_in ),
       .io_en_3( io_VwirePorts_3_3_5_en ),
       .io_en_2( io_VwirePorts_2_3_5_en ),
       .io_en_1( io_VwirePorts_1_3_5_en ),
       .io_en_0( io_VwirePorts_0_3_5_en ),
       .io_out( Vwire_164_io_out )
  );
  Vwire_2 Vwire_165(
       .io_in_3( io_VwirePorts_3_4_5_in ),
       .io_in_2( io_VwirePorts_2_4_5_in ),
       .io_in_1( io_VwirePorts_1_4_5_in ),
       .io_in_0( io_VwirePorts_0_4_5_in ),
       .io_en_3( io_VwirePorts_3_4_5_en ),
       .io_en_2( io_VwirePorts_2_4_5_en ),
       .io_en_1( io_VwirePorts_1_4_5_en ),
       .io_en_0( io_VwirePorts_0_4_5_en ),
       .io_out( Vwire_165_io_out )
  );
  Vwire_2 Vwire_166(
       .io_in_3( io_VwirePorts_3_5_5_in ),
       .io_in_2( io_VwirePorts_2_5_5_in ),
       .io_in_1( io_VwirePorts_1_5_5_in ),
       .io_in_0( io_VwirePorts_0_5_5_in ),
       .io_en_3( io_VwirePorts_3_5_5_en ),
       .io_en_2( io_VwirePorts_2_5_5_en ),
       .io_en_1( io_VwirePorts_1_5_5_en ),
       .io_en_0( io_VwirePorts_0_5_5_en ),
       .io_out( Vwire_166_io_out )
  );
  Vwire_2 Vwire_167(
       .io_in_3( io_VwirePorts_3_6_5_in ),
       .io_in_2( io_VwirePorts_2_6_5_in ),
       .io_in_1( io_VwirePorts_1_6_5_in ),
       .io_in_0( io_VwirePorts_0_6_5_in ),
       .io_en_3( io_VwirePorts_3_6_5_en ),
       .io_en_2( io_VwirePorts_2_6_5_en ),
       .io_en_1( io_VwirePorts_1_6_5_en ),
       .io_en_0( io_VwirePorts_0_6_5_en ),
       .io_out( Vwire_167_io_out )
  );
  Vwire_2 Vwire_168(
       .io_in_3( io_VwirePorts_3_7_5_in ),
       .io_in_2( io_VwirePorts_2_7_5_in ),
       .io_in_1( io_VwirePorts_1_7_5_in ),
       .io_in_0( io_VwirePorts_0_7_5_in ),
       .io_en_3( io_VwirePorts_3_7_5_en ),
       .io_en_2( io_VwirePorts_2_7_5_en ),
       .io_en_1( io_VwirePorts_1_7_5_en ),
       .io_en_0( io_VwirePorts_0_7_5_en ),
       .io_out( Vwire_168_io_out )
  );
  Vwire_2 Vwire_169(
       .io_in_3( io_VwirePorts_3_8_5_in ),
       .io_in_2( io_VwirePorts_2_8_5_in ),
       .io_in_1( io_VwirePorts_1_8_5_in ),
       .io_in_0( io_VwirePorts_0_8_5_in ),
       .io_en_3( io_VwirePorts_3_8_5_en ),
       .io_en_2( io_VwirePorts_2_8_5_en ),
       .io_en_1( io_VwirePorts_1_8_5_en ),
       .io_en_0( io_VwirePorts_0_8_5_en ),
       .io_out( Vwire_169_io_out )
  );
  Vwire_2 Vwire_170(
       .io_in_3( io_VwirePorts_3_9_5_in ),
       .io_in_2( io_VwirePorts_2_9_5_in ),
       .io_in_1( io_VwirePorts_1_9_5_in ),
       .io_in_0( io_VwirePorts_0_9_5_in ),
       .io_en_3( io_VwirePorts_3_9_5_en ),
       .io_en_2( io_VwirePorts_2_9_5_en ),
       .io_en_1( io_VwirePorts_1_9_5_en ),
       .io_en_0( io_VwirePorts_0_9_5_en ),
       .io_out( Vwire_170_io_out )
  );
  Vwire_2 Vwire_171(
       .io_in_3( io_VwirePorts_3_10_5_in ),
       .io_in_2( io_VwirePorts_2_10_5_in ),
       .io_in_1( io_VwirePorts_1_10_5_in ),
       .io_in_0( io_VwirePorts_0_10_5_in ),
       .io_en_3( io_VwirePorts_3_10_5_en ),
       .io_en_2( io_VwirePorts_2_10_5_en ),
       .io_en_1( io_VwirePorts_1_10_5_en ),
       .io_en_0( io_VwirePorts_0_10_5_en ),
       .io_out( Vwire_171_io_out )
  );
  Vwire_2 Vwire_172(
       .io_in_3( io_VwirePorts_3_11_5_in ),
       .io_in_2( io_VwirePorts_2_11_5_in ),
       .io_in_1( io_VwirePorts_1_11_5_in ),
       .io_in_0( io_VwirePorts_0_11_5_in ),
       .io_en_3( io_VwirePorts_3_11_5_en ),
       .io_en_2( io_VwirePorts_2_11_5_en ),
       .io_en_1( io_VwirePorts_1_11_5_en ),
       .io_en_0( io_VwirePorts_0_11_5_en ),
       .io_out( Vwire_172_io_out )
  );
  Vwire_2 Vwire_173(
       .io_in_3( io_VwirePorts_3_12_5_in ),
       .io_in_2( io_VwirePorts_2_12_5_in ),
       .io_in_1( io_VwirePorts_1_12_5_in ),
       .io_in_0( io_VwirePorts_0_12_5_in ),
       .io_en_3( io_VwirePorts_3_12_5_en ),
       .io_en_2( io_VwirePorts_2_12_5_en ),
       .io_en_1( io_VwirePorts_1_12_5_en ),
       .io_en_0( io_VwirePorts_0_12_5_en ),
       .io_out( Vwire_173_io_out )
  );
  Vwire_2 Vwire_174(
       .io_in_3( io_VwirePorts_3_13_5_in ),
       .io_in_2( io_VwirePorts_2_13_5_in ),
       .io_in_1( io_VwirePorts_1_13_5_in ),
       .io_in_0( io_VwirePorts_0_13_5_in ),
       .io_en_3( io_VwirePorts_3_13_5_en ),
       .io_en_2( io_VwirePorts_2_13_5_en ),
       .io_en_1( io_VwirePorts_1_13_5_en ),
       .io_en_0( io_VwirePorts_0_13_5_en ),
       .io_out( Vwire_174_io_out )
  );
  Vwire_2 Vwire_175(
       .io_in_3( io_VwirePorts_3_14_5_in ),
       .io_in_2( io_VwirePorts_2_14_5_in ),
       .io_in_1( io_VwirePorts_1_14_5_in ),
       .io_in_0( io_VwirePorts_0_14_5_in ),
       .io_en_3( io_VwirePorts_3_14_5_en ),
       .io_en_2( io_VwirePorts_2_14_5_en ),
       .io_en_1( io_VwirePorts_1_14_5_en ),
       .io_en_0( io_VwirePorts_0_14_5_en ),
       .io_out( Vwire_175_io_out )
  );
  Vwire_2 Vwire_176(
       .io_in_3( io_VwirePorts_3_15_5_in ),
       .io_in_2( io_VwirePorts_2_15_5_in ),
       .io_in_1( io_VwirePorts_1_15_5_in ),
       .io_in_0( io_VwirePorts_0_15_5_in ),
       .io_en_3( io_VwirePorts_3_15_5_en ),
       .io_en_2( io_VwirePorts_2_15_5_en ),
       .io_en_1( io_VwirePorts_1_15_5_en ),
       .io_en_0( io_VwirePorts_0_15_5_en ),
       .io_out( Vwire_176_io_out )
  );
  Vwire_2 Vwire_177(
       .io_in_3( io_VwirePorts_3_16_5_in ),
       .io_in_2( io_VwirePorts_2_16_5_in ),
       .io_in_1( io_VwirePorts_1_16_5_in ),
       .io_in_0( io_VwirePorts_0_16_5_in ),
       .io_en_3( io_VwirePorts_3_16_5_en ),
       .io_en_2( io_VwirePorts_2_16_5_en ),
       .io_en_1( io_VwirePorts_1_16_5_en ),
       .io_en_0( io_VwirePorts_0_16_5_en ),
       .io_out( Vwire_177_io_out )
  );
  Vwire_2 Vwire_178(
       .io_in_3( io_VwirePorts_3_17_5_in ),
       .io_in_2( io_VwirePorts_2_17_5_in ),
       .io_in_1( io_VwirePorts_1_17_5_in ),
       .io_in_0( io_VwirePorts_0_17_5_in ),
       .io_en_3( io_VwirePorts_3_17_5_en ),
       .io_en_2( io_VwirePorts_2_17_5_en ),
       .io_en_1( io_VwirePorts_1_17_5_en ),
       .io_en_0( io_VwirePorts_0_17_5_en ),
       .io_out( Vwire_178_io_out )
  );
  Vwire_2 Vwire_179(
       .io_in_3( io_VwirePorts_3_18_5_in ),
       .io_in_2( io_VwirePorts_2_18_5_in ),
       .io_in_1( io_VwirePorts_1_18_5_in ),
       .io_in_0( io_VwirePorts_0_18_5_in ),
       .io_en_3( io_VwirePorts_3_18_5_en ),
       .io_en_2( io_VwirePorts_2_18_5_en ),
       .io_en_1( io_VwirePorts_1_18_5_en ),
       .io_en_0( io_VwirePorts_0_18_5_en ),
       .io_out( Vwire_179_io_out )
  );
  Vwire_2 Vwire_180(
       .io_in_3( io_VwirePorts_3_19_5_in ),
       .io_in_2( io_VwirePorts_2_19_5_in ),
       .io_in_1( io_VwirePorts_1_19_5_in ),
       .io_in_0( io_VwirePorts_0_19_5_in ),
       .io_en_3( io_VwirePorts_3_19_5_en ),
       .io_en_2( io_VwirePorts_2_19_5_en ),
       .io_en_1( io_VwirePorts_1_19_5_en ),
       .io_en_0( io_VwirePorts_0_19_5_en ),
       .io_out( Vwire_180_io_out )
  );
  Vwire_2 Vwire_181(
       .io_in_3( io_VwirePorts_3_20_5_in ),
       .io_in_2( io_VwirePorts_2_20_5_in ),
       .io_in_1( io_VwirePorts_1_20_5_in ),
       .io_in_0( io_VwirePorts_0_20_5_in ),
       .io_en_3( io_VwirePorts_3_20_5_en ),
       .io_en_2( io_VwirePorts_2_20_5_en ),
       .io_en_1( io_VwirePorts_1_20_5_en ),
       .io_en_0( io_VwirePorts_0_20_5_en ),
       .io_out( Vwire_181_io_out )
  );
  Vwire_2 Vwire_182(
       .io_in_3( io_VwirePorts_3_21_5_in ),
       .io_in_2( io_VwirePorts_2_21_5_in ),
       .io_in_1( io_VwirePorts_1_21_5_in ),
       .io_in_0( io_VwirePorts_0_21_5_in ),
       .io_en_3( io_VwirePorts_3_21_5_en ),
       .io_en_2( io_VwirePorts_2_21_5_en ),
       .io_en_1( io_VwirePorts_1_21_5_en ),
       .io_en_0( io_VwirePorts_0_21_5_en ),
       .io_out( Vwire_182_io_out )
  );
  Vwire_2 Vwire_183(
       .io_in_3( io_VwirePorts_3_22_5_in ),
       .io_in_2( io_VwirePorts_2_22_5_in ),
       .io_in_1( io_VwirePorts_1_22_5_in ),
       .io_in_0( io_VwirePorts_0_22_5_in ),
       .io_en_3( io_VwirePorts_3_22_5_en ),
       .io_en_2( io_VwirePorts_2_22_5_en ),
       .io_en_1( io_VwirePorts_1_22_5_en ),
       .io_en_0( io_VwirePorts_0_22_5_en ),
       .io_out( Vwire_183_io_out )
  );
endmodule

module GarpAccel(input clk, input reset,
    input [1:0] io_mem_bus_in_23,
    input [1:0] io_mem_bus_in_22,
    input [1:0] io_mem_bus_in_21,
    input [1:0] io_mem_bus_in_20,
    input [1:0] io_mem_bus_in_19,
    input [1:0] io_mem_bus_in_18,
    input [1:0] io_mem_bus_in_17,
    input [1:0] io_mem_bus_in_16,
    input [1:0] io_mem_bus_in_15,
    input [1:0] io_mem_bus_in_14,
    input [1:0] io_mem_bus_in_13,
    input [1:0] io_mem_bus_in_12,
    input [1:0] io_mem_bus_in_11,
    input [1:0] io_mem_bus_in_10,
    input [1:0] io_mem_bus_in_9,
    input [1:0] io_mem_bus_in_8,
    input [1:0] io_mem_bus_in_7,
    input [1:0] io_mem_bus_in_6,
    input [1:0] io_mem_bus_in_5,
    input [1:0] io_mem_bus_in_4,
    input [1:0] io_mem_bus_in_3,
    input [1:0] io_mem_bus_in_2,
    input [1:0] io_mem_bus_in_1,
    input [1:0] io_mem_bus_in_0,
    output[1:0] io_mem_bus_out_23,
    output[1:0] io_mem_bus_out_22,
    output[1:0] io_mem_bus_out_21,
    output[1:0] io_mem_bus_out_20,
    output[1:0] io_mem_bus_out_19,
    output[1:0] io_mem_bus_out_18,
    output[1:0] io_mem_bus_out_17,
    output[1:0] io_mem_bus_out_16,
    output[1:0] io_mem_bus_out_15,
    output[1:0] io_mem_bus_out_14,
    output[1:0] io_mem_bus_out_13,
    output[1:0] io_mem_bus_out_12,
    output[1:0] io_mem_bus_out_11,
    output[1:0] io_mem_bus_out_10,
    output[1:0] io_mem_bus_out_9,
    output[1:0] io_mem_bus_out_8,
    output[1:0] io_mem_bus_out_7,
    output[1:0] io_mem_bus_out_6,
    output[1:0] io_mem_bus_out_5,
    output[1:0] io_mem_bus_out_4,
    output[1:0] io_mem_bus_out_3,
    output[1:0] io_mem_bus_out_2,
    output[1:0] io_mem_bus_out_1,
    output[1:0] io_mem_bus_out_0,
    input [4:0] io_addr
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire T614;
  wire T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire T684;
  wire T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire T774;
  wire T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire T790;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire T852;
  wire T853;
  wire T854;
  wire T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire T860;
  wire T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire T868;
  wire T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire T894;
  wire T895;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire T900;
  wire T901;
  wire T902;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire T916;
  wire T917;
  wire T918;
  wire T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire T924;
  wire T925;
  wire T926;
  wire T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire T932;
  wire T933;
  wire T934;
  wire T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire T940;
  wire T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire T948;
  wire T949;
  wire T950;
  wire T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire T956;
  wire T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire T964;
  wire T965;
  wire T966;
  wire T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire T972;
  wire T973;
  wire T974;
  wire T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire T980;
  wire T981;
  wire T982;
  wire T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire T988;
  wire T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire T1004;
  wire T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire T1036;
  wire T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire T1044;
  wire T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire T1052;
  wire T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire T1060;
  wire T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire T1076;
  wire T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire T1084;
  wire T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  wire T1090;
  wire T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire T1106;
  wire T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire T1113;
  wire T1114;
  wire T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire T1145;
  wire T1146;
  wire T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire T1153;
  wire T1154;
  wire T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire T1169;
  wire T1170;
  wire T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire T1185;
  wire T1186;
  wire T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire T1209;
  wire T1210;
  wire T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire T1217;
  wire T1218;
  wire T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire T1233;
  wire T1234;
  wire T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire T1257;
  wire T1258;
  wire T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire T1273;
  wire T1274;
  wire T1275;
  wire T1276;
  wire T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire T1289;
  wire T1290;
  wire T1291;
  wire T1292;
  wire T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire T1297;
  wire T1298;
  wire T1299;
  wire T1300;
  wire T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire T1305;
  wire T1306;
  wire T1307;
  wire T1308;
  wire T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire T1314;
  wire T1315;
  wire T1316;
  wire T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  wire T1324;
  wire T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire T1329;
  wire T1330;
  wire T1331;
  wire T1332;
  wire T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire T1340;
  wire T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire T1348;
  wire T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire T1353;
  wire T1354;
  wire T1355;
  wire T1356;
  wire T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire T1361;
  wire T1362;
  wire T1363;
  wire T1364;
  wire T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire T1369;
  wire T1370;
  wire T1371;
  wire T1372;
  wire T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  wire T1378;
  wire T1379;
  wire T1380;
  wire T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire T1385;
  wire T1386;
  wire T1387;
  wire T1388;
  wire T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  wire T1395;
  wire T1396;
  wire T1397;
  wire T1398;
  wire T1399;
  wire T1400;
  wire T1401;
  wire T1402;
  wire T1403;
  wire T1404;
  wire T1405;
  wire T1406;
  wire T1407;
  wire T1408;
  wire T1409;
  wire T1410;
  wire T1411;
  wire T1412;
  wire T1413;
  wire T1414;
  wire T1415;
  wire T1416;
  wire T1417;
  wire T1418;
  wire T1419;
  wire T1420;
  wire T1421;
  wire T1422;
  wire T1423;
  wire T1424;
  wire T1425;
  wire T1426;
  wire T1427;
  wire T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire T1432;
  wire T1433;
  wire T1434;
  wire T1435;
  wire T1436;
  wire T1437;
  wire T1438;
  wire T1439;
  wire T1440;
  wire T1441;
  wire T1442;
  wire T1443;
  wire T1444;
  wire T1445;
  wire T1446;
  wire T1447;
  wire T1448;
  wire T1449;
  wire T1450;
  wire T1451;
  wire T1452;
  wire T1453;
  wire T1454;
  wire T1455;
  wire T1456;
  wire T1457;
  wire T1458;
  wire T1459;
  wire T1460;
  wire T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire T1465;
  wire T1466;
  wire T1467;
  wire T1468;
  wire T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire[31:0] row_en;
  wire T1473;
  wire T1474;
  wire T1475;
  wire[1:0] T1476;
  wire[1:0] T1477;
  wire[1:0] T1478;
  wire[1:0] T1479;
  wire[1:0] T1480;
  wire[1:0] T1481;
  wire[1:0] T1482;
  wire[1:0] T1483;
  wire[1:0] T1484;
  wire[1:0] T1485;
  wire[1:0] T1486;
  wire[1:0] T1487;
  wire[1:0] T1488;
  wire[1:0] T1489;
  wire[1:0] T1490;
  wire[1:0] T1491;
  wire[1:0] T1492;
  wire[1:0] T1493;
  wire[1:0] T1494;
  wire[1:0] T1495;
  wire[1:0] T1496;
  wire[1:0] T1497;
  wire[1:0] T1498;
  wire[1:0] T1499;
  wire[1:0] T1500;
  wire[1:0] T1501;
  wire[1:0] T1502;
  wire[1:0] T1503;
  wire[1:0] T1504;
  wire[1:0] T1505;
  wire[1:0] T1506;
  wire[1:0] T1507;
  wire[1:0] T1508;
  wire[1:0] T1509;
  wire[1:0] T1510;
  wire[1:0] T1511;
  wire[1:0] T1512;
  wire[1:0] T1513;
  wire[1:0] T1514;
  wire[1:0] T1515;
  wire[1:0] T1516;
  wire[1:0] T1517;
  wire[1:0] T1518;
  wire[1:0] T1519;
  wire[1:0] T1520;
  wire[1:0] T1521;
  wire[1:0] T1522;
  wire[1:0] T1523;
  wire[1:0] T1524;
  wire[1:0] T1525;
  wire[1:0] T1526;
  wire[1:0] T1527;
  wire[1:0] T1528;
  wire[1:0] T1529;
  wire[1:0] T1530;
  wire[1:0] T1531;
  wire[1:0] T1532;
  wire[1:0] T1533;
  wire[1:0] T1534;
  wire[1:0] T1535;
  wire[31:0] ConfigAddrDecoder_io_en;
  wire[1:0] ArrayRowModule_io_V_wire_out_367;
  wire[1:0] ArrayRowModule_io_V_wire_out_366;
  wire[1:0] ArrayRowModule_io_V_wire_out_365;
  wire[1:0] ArrayRowModule_io_V_wire_out_364;
  wire[1:0] ArrayRowModule_io_V_wire_out_363;
  wire[1:0] ArrayRowModule_io_V_wire_out_362;
  wire[1:0] ArrayRowModule_io_V_wire_out_361;
  wire[1:0] ArrayRowModule_io_V_wire_out_360;
  wire[1:0] ArrayRowModule_io_V_wire_out_359;
  wire[1:0] ArrayRowModule_io_V_wire_out_358;
  wire[1:0] ArrayRowModule_io_V_wire_out_357;
  wire[1:0] ArrayRowModule_io_V_wire_out_356;
  wire[1:0] ArrayRowModule_io_V_wire_out_355;
  wire[1:0] ArrayRowModule_io_V_wire_out_354;
  wire[1:0] ArrayRowModule_io_V_wire_out_353;
  wire[1:0] ArrayRowModule_io_V_wire_out_352;
  wire[1:0] ArrayRowModule_io_V_wire_out_351;
  wire[1:0] ArrayRowModule_io_V_wire_out_350;
  wire[1:0] ArrayRowModule_io_V_wire_out_349;
  wire[1:0] ArrayRowModule_io_V_wire_out_348;
  wire[1:0] ArrayRowModule_io_V_wire_out_347;
  wire[1:0] ArrayRowModule_io_V_wire_out_346;
  wire[1:0] ArrayRowModule_io_V_wire_out_345;
  wire[1:0] ArrayRowModule_io_V_wire_out_344;
  wire[1:0] ArrayRowModule_io_V_wire_out_343;
  wire[1:0] ArrayRowModule_io_V_wire_out_342;
  wire[1:0] ArrayRowModule_io_V_wire_out_341;
  wire[1:0] ArrayRowModule_io_V_wire_out_340;
  wire[1:0] ArrayRowModule_io_V_wire_out_339;
  wire[1:0] ArrayRowModule_io_V_wire_out_338;
  wire[1:0] ArrayRowModule_io_V_wire_out_337;
  wire[1:0] ArrayRowModule_io_V_wire_out_336;
  wire[1:0] ArrayRowModule_io_V_wire_out_335;
  wire[1:0] ArrayRowModule_io_V_wire_out_334;
  wire[1:0] ArrayRowModule_io_V_wire_out_333;
  wire[1:0] ArrayRowModule_io_V_wire_out_332;
  wire[1:0] ArrayRowModule_io_V_wire_out_331;
  wire[1:0] ArrayRowModule_io_V_wire_out_330;
  wire[1:0] ArrayRowModule_io_V_wire_out_329;
  wire[1:0] ArrayRowModule_io_V_wire_out_328;
  wire[1:0] ArrayRowModule_io_V_wire_out_327;
  wire[1:0] ArrayRowModule_io_V_wire_out_326;
  wire[1:0] ArrayRowModule_io_V_wire_out_325;
  wire[1:0] ArrayRowModule_io_V_wire_out_324;
  wire[1:0] ArrayRowModule_io_V_wire_out_323;
  wire[1:0] ArrayRowModule_io_V_wire_out_322;
  wire[1:0] ArrayRowModule_io_V_wire_out_321;
  wire[1:0] ArrayRowModule_io_V_wire_out_320;
  wire[1:0] ArrayRowModule_io_V_wire_out_319;
  wire[1:0] ArrayRowModule_io_V_wire_out_318;
  wire[1:0] ArrayRowModule_io_V_wire_out_317;
  wire[1:0] ArrayRowModule_io_V_wire_out_316;
  wire[1:0] ArrayRowModule_io_V_wire_out_315;
  wire[1:0] ArrayRowModule_io_V_wire_out_314;
  wire[1:0] ArrayRowModule_io_V_wire_out_313;
  wire[1:0] ArrayRowModule_io_V_wire_out_312;
  wire[1:0] ArrayRowModule_io_V_wire_out_311;
  wire[1:0] ArrayRowModule_io_V_wire_out_310;
  wire[1:0] ArrayRowModule_io_V_wire_out_309;
  wire[1:0] ArrayRowModule_io_V_wire_out_308;
  wire[1:0] ArrayRowModule_io_V_wire_out_307;
  wire[1:0] ArrayRowModule_io_V_wire_out_306;
  wire[1:0] ArrayRowModule_io_V_wire_out_305;
  wire[1:0] ArrayRowModule_io_V_wire_out_304;
  wire[1:0] ArrayRowModule_io_V_wire_out_303;
  wire[1:0] ArrayRowModule_io_V_wire_out_302;
  wire[1:0] ArrayRowModule_io_V_wire_out_301;
  wire[1:0] ArrayRowModule_io_V_wire_out_300;
  wire[1:0] ArrayRowModule_io_V_wire_out_299;
  wire[1:0] ArrayRowModule_io_V_wire_out_298;
  wire[1:0] ArrayRowModule_io_V_wire_out_297;
  wire[1:0] ArrayRowModule_io_V_wire_out_296;
  wire[1:0] ArrayRowModule_io_V_wire_out_295;
  wire[1:0] ArrayRowModule_io_V_wire_out_294;
  wire[1:0] ArrayRowModule_io_V_wire_out_293;
  wire[1:0] ArrayRowModule_io_V_wire_out_292;
  wire[1:0] ArrayRowModule_io_V_wire_out_291;
  wire[1:0] ArrayRowModule_io_V_wire_out_290;
  wire[1:0] ArrayRowModule_io_V_wire_out_289;
  wire[1:0] ArrayRowModule_io_V_wire_out_288;
  wire[1:0] ArrayRowModule_io_V_wire_out_287;
  wire[1:0] ArrayRowModule_io_V_wire_out_286;
  wire[1:0] ArrayRowModule_io_V_wire_out_285;
  wire[1:0] ArrayRowModule_io_V_wire_out_284;
  wire[1:0] ArrayRowModule_io_V_wire_out_283;
  wire[1:0] ArrayRowModule_io_V_wire_out_282;
  wire[1:0] ArrayRowModule_io_V_wire_out_281;
  wire[1:0] ArrayRowModule_io_V_wire_out_280;
  wire[1:0] ArrayRowModule_io_V_wire_out_279;
  wire[1:0] ArrayRowModule_io_V_wire_out_278;
  wire[1:0] ArrayRowModule_io_V_wire_out_277;
  wire[1:0] ArrayRowModule_io_V_wire_out_276;
  wire[1:0] ArrayRowModule_io_V_wire_out_275;
  wire[1:0] ArrayRowModule_io_V_wire_out_274;
  wire[1:0] ArrayRowModule_io_V_wire_out_273;
  wire[1:0] ArrayRowModule_io_V_wire_out_272;
  wire[1:0] ArrayRowModule_io_V_wire_out_271;
  wire[1:0] ArrayRowModule_io_V_wire_out_270;
  wire[1:0] ArrayRowModule_io_V_wire_out_269;
  wire[1:0] ArrayRowModule_io_V_wire_out_268;
  wire[1:0] ArrayRowModule_io_V_wire_out_267;
  wire[1:0] ArrayRowModule_io_V_wire_out_266;
  wire[1:0] ArrayRowModule_io_V_wire_out_265;
  wire[1:0] ArrayRowModule_io_V_wire_out_264;
  wire[1:0] ArrayRowModule_io_V_wire_out_263;
  wire[1:0] ArrayRowModule_io_V_wire_out_262;
  wire[1:0] ArrayRowModule_io_V_wire_out_261;
  wire[1:0] ArrayRowModule_io_V_wire_out_260;
  wire[1:0] ArrayRowModule_io_V_wire_out_259;
  wire[1:0] ArrayRowModule_io_V_wire_out_258;
  wire[1:0] ArrayRowModule_io_V_wire_out_257;
  wire[1:0] ArrayRowModule_io_V_wire_out_256;
  wire[1:0] ArrayRowModule_io_V_wire_out_255;
  wire[1:0] ArrayRowModule_io_V_wire_out_254;
  wire[1:0] ArrayRowModule_io_V_wire_out_253;
  wire[1:0] ArrayRowModule_io_V_wire_out_252;
  wire[1:0] ArrayRowModule_io_V_wire_out_251;
  wire[1:0] ArrayRowModule_io_V_wire_out_250;
  wire[1:0] ArrayRowModule_io_V_wire_out_249;
  wire[1:0] ArrayRowModule_io_V_wire_out_248;
  wire[1:0] ArrayRowModule_io_V_wire_out_247;
  wire[1:0] ArrayRowModule_io_V_wire_out_246;
  wire[1:0] ArrayRowModule_io_V_wire_out_245;
  wire[1:0] ArrayRowModule_io_V_wire_out_244;
  wire[1:0] ArrayRowModule_io_V_wire_out_243;
  wire[1:0] ArrayRowModule_io_V_wire_out_242;
  wire[1:0] ArrayRowModule_io_V_wire_out_241;
  wire[1:0] ArrayRowModule_io_V_wire_out_240;
  wire[1:0] ArrayRowModule_io_V_wire_out_239;
  wire[1:0] ArrayRowModule_io_V_wire_out_238;
  wire[1:0] ArrayRowModule_io_V_wire_out_237;
  wire[1:0] ArrayRowModule_io_V_wire_out_236;
  wire[1:0] ArrayRowModule_io_V_wire_out_235;
  wire[1:0] ArrayRowModule_io_V_wire_out_234;
  wire[1:0] ArrayRowModule_io_V_wire_out_233;
  wire[1:0] ArrayRowModule_io_V_wire_out_232;
  wire[1:0] ArrayRowModule_io_V_wire_out_231;
  wire[1:0] ArrayRowModule_io_V_wire_out_230;
  wire[1:0] ArrayRowModule_io_V_wire_out_229;
  wire[1:0] ArrayRowModule_io_V_wire_out_228;
  wire[1:0] ArrayRowModule_io_V_wire_out_227;
  wire[1:0] ArrayRowModule_io_V_wire_out_226;
  wire[1:0] ArrayRowModule_io_V_wire_out_225;
  wire[1:0] ArrayRowModule_io_V_wire_out_224;
  wire[1:0] ArrayRowModule_io_V_wire_out_223;
  wire[1:0] ArrayRowModule_io_V_wire_out_222;
  wire[1:0] ArrayRowModule_io_V_wire_out_221;
  wire[1:0] ArrayRowModule_io_V_wire_out_220;
  wire[1:0] ArrayRowModule_io_V_wire_out_219;
  wire[1:0] ArrayRowModule_io_V_wire_out_218;
  wire[1:0] ArrayRowModule_io_V_wire_out_217;
  wire[1:0] ArrayRowModule_io_V_wire_out_216;
  wire[1:0] ArrayRowModule_io_V_wire_out_215;
  wire[1:0] ArrayRowModule_io_V_wire_out_214;
  wire[1:0] ArrayRowModule_io_V_wire_out_213;
  wire[1:0] ArrayRowModule_io_V_wire_out_212;
  wire[1:0] ArrayRowModule_io_V_wire_out_211;
  wire[1:0] ArrayRowModule_io_V_wire_out_210;
  wire[1:0] ArrayRowModule_io_V_wire_out_209;
  wire[1:0] ArrayRowModule_io_V_wire_out_208;
  wire[1:0] ArrayRowModule_io_V_wire_out_207;
  wire[1:0] ArrayRowModule_io_V_wire_out_206;
  wire[1:0] ArrayRowModule_io_V_wire_out_205;
  wire[1:0] ArrayRowModule_io_V_wire_out_204;
  wire[1:0] ArrayRowModule_io_V_wire_out_203;
  wire[1:0] ArrayRowModule_io_V_wire_out_202;
  wire[1:0] ArrayRowModule_io_V_wire_out_201;
  wire[1:0] ArrayRowModule_io_V_wire_out_200;
  wire[1:0] ArrayRowModule_io_V_wire_out_199;
  wire[1:0] ArrayRowModule_io_V_wire_out_198;
  wire[1:0] ArrayRowModule_io_V_wire_out_197;
  wire[1:0] ArrayRowModule_io_V_wire_out_196;
  wire[1:0] ArrayRowModule_io_V_wire_out_195;
  wire[1:0] ArrayRowModule_io_V_wire_out_194;
  wire[1:0] ArrayRowModule_io_V_wire_out_193;
  wire[1:0] ArrayRowModule_io_V_wire_out_192;
  wire[1:0] ArrayRowModule_io_V_wire_out_191;
  wire[1:0] ArrayRowModule_io_V_wire_out_190;
  wire[1:0] ArrayRowModule_io_V_wire_out_189;
  wire[1:0] ArrayRowModule_io_V_wire_out_188;
  wire[1:0] ArrayRowModule_io_V_wire_out_187;
  wire[1:0] ArrayRowModule_io_V_wire_out_186;
  wire[1:0] ArrayRowModule_io_V_wire_out_185;
  wire[1:0] ArrayRowModule_io_V_wire_out_184;
  wire[1:0] ArrayRowModule_io_V_wire_out_183;
  wire[1:0] ArrayRowModule_io_V_wire_out_182;
  wire[1:0] ArrayRowModule_io_V_wire_out_181;
  wire[1:0] ArrayRowModule_io_V_wire_out_180;
  wire[1:0] ArrayRowModule_io_V_wire_out_179;
  wire[1:0] ArrayRowModule_io_V_wire_out_178;
  wire[1:0] ArrayRowModule_io_V_wire_out_177;
  wire[1:0] ArrayRowModule_io_V_wire_out_176;
  wire[1:0] ArrayRowModule_io_V_wire_out_175;
  wire[1:0] ArrayRowModule_io_V_wire_out_174;
  wire[1:0] ArrayRowModule_io_V_wire_out_173;
  wire[1:0] ArrayRowModule_io_V_wire_out_172;
  wire[1:0] ArrayRowModule_io_V_wire_out_171;
  wire[1:0] ArrayRowModule_io_V_wire_out_170;
  wire[1:0] ArrayRowModule_io_V_wire_out_169;
  wire[1:0] ArrayRowModule_io_V_wire_out_168;
  wire[1:0] ArrayRowModule_io_V_wire_out_167;
  wire[1:0] ArrayRowModule_io_V_wire_out_166;
  wire[1:0] ArrayRowModule_io_V_wire_out_165;
  wire[1:0] ArrayRowModule_io_V_wire_out_164;
  wire[1:0] ArrayRowModule_io_V_wire_out_163;
  wire[1:0] ArrayRowModule_io_V_wire_out_162;
  wire[1:0] ArrayRowModule_io_V_wire_out_161;
  wire[1:0] ArrayRowModule_io_V_wire_out_160;
  wire[1:0] ArrayRowModule_io_V_wire_out_159;
  wire[1:0] ArrayRowModule_io_V_wire_out_158;
  wire[1:0] ArrayRowModule_io_V_wire_out_157;
  wire[1:0] ArrayRowModule_io_V_wire_out_156;
  wire[1:0] ArrayRowModule_io_V_wire_out_155;
  wire[1:0] ArrayRowModule_io_V_wire_out_154;
  wire[1:0] ArrayRowModule_io_V_wire_out_153;
  wire[1:0] ArrayRowModule_io_V_wire_out_152;
  wire[1:0] ArrayRowModule_io_V_wire_out_151;
  wire[1:0] ArrayRowModule_io_V_wire_out_150;
  wire[1:0] ArrayRowModule_io_V_wire_out_149;
  wire[1:0] ArrayRowModule_io_V_wire_out_148;
  wire[1:0] ArrayRowModule_io_V_wire_out_147;
  wire[1:0] ArrayRowModule_io_V_wire_out_146;
  wire[1:0] ArrayRowModule_io_V_wire_out_145;
  wire[1:0] ArrayRowModule_io_V_wire_out_144;
  wire[1:0] ArrayRowModule_io_V_wire_out_143;
  wire[1:0] ArrayRowModule_io_V_wire_out_142;
  wire[1:0] ArrayRowModule_io_V_wire_out_141;
  wire[1:0] ArrayRowModule_io_V_wire_out_140;
  wire[1:0] ArrayRowModule_io_V_wire_out_139;
  wire[1:0] ArrayRowModule_io_V_wire_out_138;
  wire[1:0] ArrayRowModule_io_V_wire_out_137;
  wire[1:0] ArrayRowModule_io_V_wire_out_136;
  wire[1:0] ArrayRowModule_io_V_wire_out_135;
  wire[1:0] ArrayRowModule_io_V_wire_out_134;
  wire[1:0] ArrayRowModule_io_V_wire_out_133;
  wire[1:0] ArrayRowModule_io_V_wire_out_132;
  wire[1:0] ArrayRowModule_io_V_wire_out_131;
  wire[1:0] ArrayRowModule_io_V_wire_out_130;
  wire[1:0] ArrayRowModule_io_V_wire_out_129;
  wire[1:0] ArrayRowModule_io_V_wire_out_128;
  wire[1:0] ArrayRowModule_io_V_wire_out_127;
  wire[1:0] ArrayRowModule_io_V_wire_out_126;
  wire[1:0] ArrayRowModule_io_V_wire_out_125;
  wire[1:0] ArrayRowModule_io_V_wire_out_124;
  wire[1:0] ArrayRowModule_io_V_wire_out_123;
  wire[1:0] ArrayRowModule_io_V_wire_out_122;
  wire[1:0] ArrayRowModule_io_V_wire_out_121;
  wire[1:0] ArrayRowModule_io_V_wire_out_120;
  wire[1:0] ArrayRowModule_io_V_wire_out_119;
  wire[1:0] ArrayRowModule_io_V_wire_out_118;
  wire[1:0] ArrayRowModule_io_V_wire_out_117;
  wire[1:0] ArrayRowModule_io_V_wire_out_116;
  wire[1:0] ArrayRowModule_io_V_wire_out_115;
  wire[1:0] ArrayRowModule_io_V_wire_out_114;
  wire[1:0] ArrayRowModule_io_V_wire_out_113;
  wire[1:0] ArrayRowModule_io_V_wire_out_112;
  wire[1:0] ArrayRowModule_io_V_wire_out_111;
  wire[1:0] ArrayRowModule_io_V_wire_out_110;
  wire[1:0] ArrayRowModule_io_V_wire_out_109;
  wire[1:0] ArrayRowModule_io_V_wire_out_108;
  wire[1:0] ArrayRowModule_io_V_wire_out_107;
  wire[1:0] ArrayRowModule_io_V_wire_out_106;
  wire[1:0] ArrayRowModule_io_V_wire_out_105;
  wire[1:0] ArrayRowModule_io_V_wire_out_104;
  wire[1:0] ArrayRowModule_io_V_wire_out_103;
  wire[1:0] ArrayRowModule_io_V_wire_out_102;
  wire[1:0] ArrayRowModule_io_V_wire_out_101;
  wire[1:0] ArrayRowModule_io_V_wire_out_100;
  wire[1:0] ArrayRowModule_io_V_wire_out_99;
  wire[1:0] ArrayRowModule_io_V_wire_out_98;
  wire[1:0] ArrayRowModule_io_V_wire_out_97;
  wire[1:0] ArrayRowModule_io_V_wire_out_96;
  wire[1:0] ArrayRowModule_io_V_wire_out_95;
  wire[1:0] ArrayRowModule_io_V_wire_out_94;
  wire[1:0] ArrayRowModule_io_V_wire_out_93;
  wire[1:0] ArrayRowModule_io_V_wire_out_92;
  wire[1:0] ArrayRowModule_io_V_wire_out_91;
  wire[1:0] ArrayRowModule_io_V_wire_out_90;
  wire[1:0] ArrayRowModule_io_V_wire_out_89;
  wire[1:0] ArrayRowModule_io_V_wire_out_88;
  wire[1:0] ArrayRowModule_io_V_wire_out_87;
  wire[1:0] ArrayRowModule_io_V_wire_out_86;
  wire[1:0] ArrayRowModule_io_V_wire_out_85;
  wire[1:0] ArrayRowModule_io_V_wire_out_84;
  wire[1:0] ArrayRowModule_io_V_wire_out_83;
  wire[1:0] ArrayRowModule_io_V_wire_out_82;
  wire[1:0] ArrayRowModule_io_V_wire_out_81;
  wire[1:0] ArrayRowModule_io_V_wire_out_80;
  wire[1:0] ArrayRowModule_io_V_wire_out_79;
  wire[1:0] ArrayRowModule_io_V_wire_out_78;
  wire[1:0] ArrayRowModule_io_V_wire_out_77;
  wire[1:0] ArrayRowModule_io_V_wire_out_76;
  wire[1:0] ArrayRowModule_io_V_wire_out_75;
  wire[1:0] ArrayRowModule_io_V_wire_out_74;
  wire[1:0] ArrayRowModule_io_V_wire_out_73;
  wire[1:0] ArrayRowModule_io_V_wire_out_72;
  wire[1:0] ArrayRowModule_io_V_wire_out_71;
  wire[1:0] ArrayRowModule_io_V_wire_out_70;
  wire[1:0] ArrayRowModule_io_V_wire_out_69;
  wire[1:0] ArrayRowModule_io_V_wire_out_68;
  wire[1:0] ArrayRowModule_io_V_wire_out_67;
  wire[1:0] ArrayRowModule_io_V_wire_out_66;
  wire[1:0] ArrayRowModule_io_V_wire_out_65;
  wire[1:0] ArrayRowModule_io_V_wire_out_64;
  wire[1:0] ArrayRowModule_io_V_wire_out_63;
  wire[1:0] ArrayRowModule_io_V_wire_out_62;
  wire[1:0] ArrayRowModule_io_V_wire_out_61;
  wire[1:0] ArrayRowModule_io_V_wire_out_60;
  wire[1:0] ArrayRowModule_io_V_wire_out_59;
  wire[1:0] ArrayRowModule_io_V_wire_out_58;
  wire[1:0] ArrayRowModule_io_V_wire_out_57;
  wire[1:0] ArrayRowModule_io_V_wire_out_56;
  wire[1:0] ArrayRowModule_io_V_wire_out_55;
  wire[1:0] ArrayRowModule_io_V_wire_out_54;
  wire[1:0] ArrayRowModule_io_V_wire_out_53;
  wire[1:0] ArrayRowModule_io_V_wire_out_52;
  wire[1:0] ArrayRowModule_io_V_wire_out_51;
  wire[1:0] ArrayRowModule_io_V_wire_out_50;
  wire[1:0] ArrayRowModule_io_V_wire_out_49;
  wire[1:0] ArrayRowModule_io_V_wire_out_48;
  wire[1:0] ArrayRowModule_io_V_wire_out_47;
  wire[1:0] ArrayRowModule_io_V_wire_out_46;
  wire[1:0] ArrayRowModule_io_V_wire_out_45;
  wire[1:0] ArrayRowModule_io_V_wire_out_44;
  wire[1:0] ArrayRowModule_io_V_wire_out_43;
  wire[1:0] ArrayRowModule_io_V_wire_out_42;
  wire[1:0] ArrayRowModule_io_V_wire_out_41;
  wire[1:0] ArrayRowModule_io_V_wire_out_40;
  wire[1:0] ArrayRowModule_io_V_wire_out_39;
  wire[1:0] ArrayRowModule_io_V_wire_out_38;
  wire[1:0] ArrayRowModule_io_V_wire_out_37;
  wire[1:0] ArrayRowModule_io_V_wire_out_36;
  wire[1:0] ArrayRowModule_io_V_wire_out_35;
  wire[1:0] ArrayRowModule_io_V_wire_out_34;
  wire[1:0] ArrayRowModule_io_V_wire_out_33;
  wire[1:0] ArrayRowModule_io_V_wire_out_32;
  wire[1:0] ArrayRowModule_io_V_wire_out_31;
  wire[1:0] ArrayRowModule_io_V_wire_out_30;
  wire[1:0] ArrayRowModule_io_V_wire_out_29;
  wire[1:0] ArrayRowModule_io_V_wire_out_28;
  wire[1:0] ArrayRowModule_io_V_wire_out_27;
  wire[1:0] ArrayRowModule_io_V_wire_out_26;
  wire[1:0] ArrayRowModule_io_V_wire_out_25;
  wire[1:0] ArrayRowModule_io_V_wire_out_24;
  wire[1:0] ArrayRowModule_io_V_wire_out_23;
  wire[1:0] ArrayRowModule_io_V_wire_out_22;
  wire[1:0] ArrayRowModule_io_V_wire_out_21;
  wire[1:0] ArrayRowModule_io_V_wire_out_20;
  wire[1:0] ArrayRowModule_io_V_wire_out_19;
  wire[1:0] ArrayRowModule_io_V_wire_out_18;
  wire[1:0] ArrayRowModule_io_V_wire_out_17;
  wire[1:0] ArrayRowModule_io_V_wire_out_16;
  wire[1:0] ArrayRowModule_io_V_wire_out_15;
  wire[1:0] ArrayRowModule_io_V_wire_out_14;
  wire[1:0] ArrayRowModule_io_V_wire_out_13;
  wire[1:0] ArrayRowModule_io_V_wire_out_12;
  wire[1:0] ArrayRowModule_io_V_wire_out_11;
  wire[1:0] ArrayRowModule_io_V_wire_out_10;
  wire[1:0] ArrayRowModule_io_V_wire_out_9;
  wire[1:0] ArrayRowModule_io_V_wire_out_8;
  wire[1:0] ArrayRowModule_io_V_wire_out_7;
  wire[1:0] ArrayRowModule_io_V_wire_out_6;
  wire[1:0] ArrayRowModule_io_V_wire_out_5;
  wire[1:0] ArrayRowModule_io_V_wire_out_4;
  wire[1:0] ArrayRowModule_io_V_wire_out_3;
  wire[1:0] ArrayRowModule_io_V_wire_out_2;
  wire[1:0] ArrayRowModule_io_V_wire_out_1;
  wire[1:0] ArrayRowModule_io_V_wire_out_0;
  wire[15:0] ArrayRowModule_io_V_wire_en_22;
  wire[15:0] ArrayRowModule_io_V_wire_en_21;
  wire[15:0] ArrayRowModule_io_V_wire_en_20;
  wire[15:0] ArrayRowModule_io_V_wire_en_19;
  wire[15:0] ArrayRowModule_io_V_wire_en_18;
  wire[15:0] ArrayRowModule_io_V_wire_en_17;
  wire[15:0] ArrayRowModule_io_V_wire_en_16;
  wire[15:0] ArrayRowModule_io_V_wire_en_15;
  wire[15:0] ArrayRowModule_io_V_wire_en_14;
  wire[15:0] ArrayRowModule_io_V_wire_en_13;
  wire[15:0] ArrayRowModule_io_V_wire_en_12;
  wire[15:0] ArrayRowModule_io_V_wire_en_11;
  wire[15:0] ArrayRowModule_io_V_wire_en_10;
  wire[15:0] ArrayRowModule_io_V_wire_en_9;
  wire[15:0] ArrayRowModule_io_V_wire_en_8;
  wire[15:0] ArrayRowModule_io_V_wire_en_7;
  wire[15:0] ArrayRowModule_io_V_wire_en_6;
  wire[15:0] ArrayRowModule_io_V_wire_en_5;
  wire[15:0] ArrayRowModule_io_V_wire_en_4;
  wire[15:0] ArrayRowModule_io_V_wire_en_3;
  wire[15:0] ArrayRowModule_io_V_wire_en_2;
  wire[15:0] ArrayRowModule_io_V_wire_en_1;
  wire[15:0] ArrayRowModule_io_V_wire_en_0;
  wire[1:0] ArrayRowModule_io_H_out_22;
  wire[1:0] ArrayRowModule_io_H_out_21;
  wire[1:0] ArrayRowModule_io_H_out_20;
  wire[1:0] ArrayRowModule_io_H_out_19;
  wire[1:0] ArrayRowModule_io_H_out_18;
  wire[1:0] ArrayRowModule_io_H_out_17;
  wire[1:0] ArrayRowModule_io_H_out_16;
  wire[1:0] ArrayRowModule_io_H_out_15;
  wire[1:0] ArrayRowModule_io_H_out_14;
  wire[1:0] ArrayRowModule_io_H_out_13;
  wire[1:0] ArrayRowModule_io_H_out_12;
  wire[1:0] ArrayRowModule_io_H_out_11;
  wire[1:0] ArrayRowModule_io_H_out_10;
  wire[1:0] ArrayRowModule_io_H_out_9;
  wire[1:0] ArrayRowModule_io_H_out_8;
  wire[1:0] ArrayRowModule_io_H_out_7;
  wire[1:0] ArrayRowModule_io_H_out_6;
  wire[1:0] ArrayRowModule_io_H_out_5;
  wire[1:0] ArrayRowModule_io_H_out_4;
  wire[1:0] ArrayRowModule_io_H_out_3;
  wire[1:0] ArrayRowModule_io_H_out_2;
  wire[1:0] ArrayRowModule_io_H_out_1;
  wire[1:0] ArrayRowModule_io_H_out_0;
  wire[1:0] ArrayRowModule_io_G_wire_below_3;
  wire[1:0] ArrayRowModule_io_G_wire_below_2;
  wire[1:0] ArrayRowModule_io_G_wire_below_1;
  wire[1:0] ArrayRowModule_io_G_wire_below_0;
  wire[1:0] ArrayRowModule_io_H_wire_below_32;
  wire[1:0] ArrayRowModule_io_H_wire_below_31;
  wire[1:0] ArrayRowModule_io_H_wire_below_30;
  wire[1:0] ArrayRowModule_io_H_wire_below_29;
  wire[1:0] ArrayRowModule_io_H_wire_below_28;
  wire[1:0] ArrayRowModule_io_H_wire_below_27;
  wire[1:0] ArrayRowModule_io_H_wire_below_26;
  wire[1:0] ArrayRowModule_io_H_wire_below_25;
  wire[1:0] ArrayRowModule_io_H_wire_below_24;
  wire[1:0] ArrayRowModule_io_H_wire_below_23;
  wire[1:0] ArrayRowModule_io_H_wire_below_22;
  wire[1:0] ArrayRowModule_io_H_wire_below_21;
  wire[1:0] ArrayRowModule_io_H_wire_below_20;
  wire[1:0] ArrayRowModule_io_H_wire_below_19;
  wire[1:0] ArrayRowModule_io_H_wire_below_18;
  wire[1:0] ArrayRowModule_io_H_wire_below_17;
  wire[1:0] ArrayRowModule_io_H_wire_below_16;
  wire[1:0] ArrayRowModule_io_H_wire_below_15;
  wire[1:0] ArrayRowModule_io_H_wire_below_14;
  wire[1:0] ArrayRowModule_io_H_wire_below_13;
  wire[1:0] ArrayRowModule_io_H_wire_below_12;
  wire[1:0] ArrayRowModule_io_H_wire_below_11;
  wire[1:0] ArrayRowModule_io_H_wire_below_10;
  wire[1:0] ArrayRowModule_io_H_wire_below_9;
  wire[1:0] ArrayRowModule_io_H_wire_below_8;
  wire[1:0] ArrayRowModule_io_H_wire_below_7;
  wire[1:0] ArrayRowModule_io_H_wire_below_6;
  wire[1:0] ArrayRowModule_io_H_wire_below_5;
  wire[1:0] ArrayRowModule_io_H_wire_below_4;
  wire[1:0] ArrayRowModule_io_H_wire_below_3;
  wire[1:0] ArrayRowModule_io_H_wire_below_2;
  wire[1:0] ArrayRowModule_io_H_wire_below_1;
  wire[1:0] ArrayRowModule_io_H_wire_below_0;
  wire[1:0] ArrayRowModule_io_mem_bus_out_23;
  wire[1:0] ArrayRowModule_io_mem_bus_out_22;
  wire[1:0] ArrayRowModule_io_mem_bus_out_21;
  wire[1:0] ArrayRowModule_io_mem_bus_out_20;
  wire[1:0] ArrayRowModule_io_mem_bus_out_19;
  wire[1:0] ArrayRowModule_io_mem_bus_out_18;
  wire[1:0] ArrayRowModule_io_mem_bus_out_17;
  wire[1:0] ArrayRowModule_io_mem_bus_out_16;
  wire[1:0] ArrayRowModule_io_mem_bus_out_15;
  wire[1:0] ArrayRowModule_io_mem_bus_out_14;
  wire[1:0] ArrayRowModule_io_mem_bus_out_13;
  wire[1:0] ArrayRowModule_io_mem_bus_out_12;
  wire[1:0] ArrayRowModule_io_mem_bus_out_11;
  wire[1:0] ArrayRowModule_io_mem_bus_out_10;
  wire[1:0] ArrayRowModule_io_mem_bus_out_9;
  wire[1:0] ArrayRowModule_io_mem_bus_out_8;
  wire[1:0] ArrayRowModule_io_mem_bus_out_7;
  wire[1:0] ArrayRowModule_io_mem_bus_out_6;
  wire[1:0] ArrayRowModule_io_mem_bus_out_5;
  wire[1:0] ArrayRowModule_io_mem_bus_out_4;
  wire[1:0] ArrayRowModule_io_mem_bus_out_3;
  wire[1:0] ArrayRowModule_io_mem_bus_out_2;
  wire[1:0] ArrayRowModule_io_mem_bus_out_1;
  wire[1:0] ArrayRowModule_io_mem_bus_out_0;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_367;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_366;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_365;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_364;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_363;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_362;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_361;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_360;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_359;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_358;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_357;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_356;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_355;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_354;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_353;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_352;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_351;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_350;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_349;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_348;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_347;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_346;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_345;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_344;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_343;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_342;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_341;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_340;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_339;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_338;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_337;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_336;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_335;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_334;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_333;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_332;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_331;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_330;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_329;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_328;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_327;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_326;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_325;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_324;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_323;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_322;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_321;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_320;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_319;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_318;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_317;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_316;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_315;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_314;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_313;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_312;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_311;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_310;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_309;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_308;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_307;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_306;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_305;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_304;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_303;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_302;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_301;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_300;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_299;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_298;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_297;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_296;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_295;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_294;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_293;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_292;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_291;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_290;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_289;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_288;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_287;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_286;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_285;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_284;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_283;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_282;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_281;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_280;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_279;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_278;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_277;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_276;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_275;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_274;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_273;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_272;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_271;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_270;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_269;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_268;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_267;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_266;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_265;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_264;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_263;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_262;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_261;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_260;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_259;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_258;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_257;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_256;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_255;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_254;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_253;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_252;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_251;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_250;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_249;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_248;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_247;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_246;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_245;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_244;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_243;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_242;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_241;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_240;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_239;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_238;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_237;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_236;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_235;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_234;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_233;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_232;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_231;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_230;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_229;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_228;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_227;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_226;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_225;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_224;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_223;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_222;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_221;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_220;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_219;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_218;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_217;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_216;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_215;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_214;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_213;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_212;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_211;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_210;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_209;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_208;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_207;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_206;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_205;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_204;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_203;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_202;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_201;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_200;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_199;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_198;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_197;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_196;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_195;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_194;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_193;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_192;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_191;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_190;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_189;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_188;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_187;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_186;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_185;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_184;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_183;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_182;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_181;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_180;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_179;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_178;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_177;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_176;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_175;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_174;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_173;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_172;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_171;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_170;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_169;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_168;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_167;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_166;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_165;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_164;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_163;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_162;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_161;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_160;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_159;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_158;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_157;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_156;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_155;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_154;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_153;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_152;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_151;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_150;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_149;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_148;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_147;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_146;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_145;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_144;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_143;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_142;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_141;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_140;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_139;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_138;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_137;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_136;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_135;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_134;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_133;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_132;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_131;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_130;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_129;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_128;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_127;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_126;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_125;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_124;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_123;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_122;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_121;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_120;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_119;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_118;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_117;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_116;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_115;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_114;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_113;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_112;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_111;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_110;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_109;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_108;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_107;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_106;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_105;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_104;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_103;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_102;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_101;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_100;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_99;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_98;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_97;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_96;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_95;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_94;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_93;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_92;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_91;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_90;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_89;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_88;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_87;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_86;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_85;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_84;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_83;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_82;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_81;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_80;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_79;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_78;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_77;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_76;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_75;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_74;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_73;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_72;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_71;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_70;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_69;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_68;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_67;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_66;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_65;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_64;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_63;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_62;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_61;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_60;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_59;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_58;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_57;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_56;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_55;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_54;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_53;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_52;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_51;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_50;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_49;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_48;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_47;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_46;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_45;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_44;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_43;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_42;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_41;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_40;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_39;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_38;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_37;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_36;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_35;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_34;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_33;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_32;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_31;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_30;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_29;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_28;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_27;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_26;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_25;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_24;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_23;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_22;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_21;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_20;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_19;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_18;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_17;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_16;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_15;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_14;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_13;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_12;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_11;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_10;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_9;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_8;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_7;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_6;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_5;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_4;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_3;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_2;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_1;
  wire[1:0] ArrayRowModule_1_io_V_wire_out_0;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_22;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_21;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_20;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_19;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_18;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_17;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_16;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_15;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_14;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_13;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_12;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_11;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_10;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_9;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_8;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_7;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_6;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_5;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_4;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_3;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_2;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_1;
  wire[15:0] ArrayRowModule_1_io_V_wire_en_0;
  wire[1:0] ArrayRowModule_1_io_H_out_22;
  wire[1:0] ArrayRowModule_1_io_H_out_21;
  wire[1:0] ArrayRowModule_1_io_H_out_20;
  wire[1:0] ArrayRowModule_1_io_H_out_19;
  wire[1:0] ArrayRowModule_1_io_H_out_18;
  wire[1:0] ArrayRowModule_1_io_H_out_17;
  wire[1:0] ArrayRowModule_1_io_H_out_16;
  wire[1:0] ArrayRowModule_1_io_H_out_15;
  wire[1:0] ArrayRowModule_1_io_H_out_14;
  wire[1:0] ArrayRowModule_1_io_H_out_13;
  wire[1:0] ArrayRowModule_1_io_H_out_12;
  wire[1:0] ArrayRowModule_1_io_H_out_11;
  wire[1:0] ArrayRowModule_1_io_H_out_10;
  wire[1:0] ArrayRowModule_1_io_H_out_9;
  wire[1:0] ArrayRowModule_1_io_H_out_8;
  wire[1:0] ArrayRowModule_1_io_H_out_7;
  wire[1:0] ArrayRowModule_1_io_H_out_6;
  wire[1:0] ArrayRowModule_1_io_H_out_5;
  wire[1:0] ArrayRowModule_1_io_H_out_4;
  wire[1:0] ArrayRowModule_1_io_H_out_3;
  wire[1:0] ArrayRowModule_1_io_H_out_2;
  wire[1:0] ArrayRowModule_1_io_H_out_1;
  wire[1:0] ArrayRowModule_1_io_H_out_0;
  wire[1:0] ArrayRowModule_1_io_G_wire_below_3;
  wire[1:0] ArrayRowModule_1_io_G_wire_below_2;
  wire[1:0] ArrayRowModule_1_io_G_wire_below_1;
  wire[1:0] ArrayRowModule_1_io_G_wire_below_0;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_32;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_31;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_30;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_29;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_28;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_27;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_26;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_25;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_24;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_23;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_22;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_21;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_20;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_19;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_18;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_17;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_16;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_15;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_14;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_13;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_12;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_11;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_10;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_9;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_8;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_7;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_6;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_5;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_4;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_3;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_2;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_1;
  wire[1:0] ArrayRowModule_1_io_H_wire_below_0;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_23;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_22;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_21;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_20;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_19;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_18;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_17;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_16;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_15;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_14;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_13;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_12;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_11;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_10;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_9;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_8;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_7;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_6;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_5;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_4;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_3;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_2;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_1;
  wire[1:0] ArrayRowModule_1_io_mem_bus_out_0;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_367;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_366;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_365;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_364;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_363;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_362;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_361;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_360;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_359;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_358;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_357;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_356;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_355;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_354;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_353;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_352;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_351;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_350;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_349;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_348;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_347;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_346;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_345;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_344;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_343;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_342;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_341;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_340;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_339;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_338;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_337;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_336;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_335;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_334;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_333;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_332;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_331;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_330;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_329;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_328;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_327;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_326;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_325;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_324;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_323;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_322;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_321;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_320;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_319;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_318;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_317;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_316;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_315;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_314;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_313;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_312;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_311;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_310;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_309;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_308;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_307;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_306;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_305;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_304;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_303;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_302;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_301;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_300;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_299;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_298;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_297;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_296;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_295;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_294;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_293;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_292;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_291;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_290;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_289;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_288;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_287;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_286;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_285;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_284;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_283;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_282;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_281;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_280;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_279;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_278;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_277;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_276;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_275;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_274;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_273;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_272;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_271;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_270;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_269;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_268;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_267;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_266;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_265;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_264;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_263;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_262;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_261;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_260;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_259;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_258;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_257;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_256;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_255;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_254;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_253;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_252;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_251;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_250;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_249;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_248;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_247;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_246;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_245;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_244;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_243;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_242;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_241;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_240;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_239;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_238;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_237;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_236;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_235;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_234;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_233;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_232;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_231;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_230;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_229;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_228;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_227;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_226;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_225;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_224;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_223;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_222;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_221;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_220;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_219;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_218;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_217;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_216;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_215;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_214;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_213;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_212;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_211;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_210;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_209;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_208;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_207;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_206;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_205;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_204;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_203;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_202;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_201;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_200;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_199;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_198;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_197;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_196;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_195;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_194;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_193;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_192;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_191;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_190;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_189;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_188;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_187;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_186;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_185;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_184;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_183;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_182;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_181;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_180;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_179;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_178;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_177;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_176;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_175;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_174;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_173;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_172;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_171;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_170;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_169;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_168;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_167;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_166;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_165;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_164;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_163;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_162;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_161;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_160;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_159;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_158;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_157;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_156;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_155;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_154;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_153;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_152;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_151;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_150;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_149;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_148;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_147;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_146;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_145;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_144;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_143;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_142;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_141;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_140;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_139;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_138;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_137;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_136;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_135;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_134;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_133;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_132;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_131;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_130;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_129;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_128;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_127;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_126;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_125;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_124;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_123;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_122;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_121;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_120;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_119;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_118;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_117;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_116;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_115;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_114;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_113;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_112;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_111;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_110;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_109;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_108;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_107;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_106;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_105;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_104;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_103;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_102;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_101;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_100;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_99;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_98;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_97;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_96;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_95;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_94;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_93;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_92;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_91;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_90;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_89;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_88;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_87;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_86;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_85;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_84;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_83;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_82;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_81;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_80;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_79;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_78;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_77;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_76;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_75;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_74;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_73;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_72;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_71;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_70;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_69;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_68;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_67;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_66;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_65;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_64;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_63;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_62;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_61;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_60;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_59;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_58;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_57;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_56;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_55;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_54;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_53;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_52;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_51;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_50;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_49;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_48;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_47;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_46;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_45;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_44;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_43;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_42;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_41;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_40;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_39;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_38;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_37;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_36;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_35;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_34;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_33;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_32;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_31;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_30;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_29;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_28;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_27;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_26;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_25;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_24;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_23;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_22;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_21;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_20;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_19;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_18;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_17;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_16;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_15;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_14;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_13;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_12;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_11;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_10;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_9;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_8;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_7;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_6;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_5;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_4;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_3;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_2;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_1;
  wire[1:0] ArrayRowModule_2_io_V_wire_out_0;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_22;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_21;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_20;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_19;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_18;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_17;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_16;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_15;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_14;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_13;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_12;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_11;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_10;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_9;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_8;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_7;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_6;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_5;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_4;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_3;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_2;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_1;
  wire[15:0] ArrayRowModule_2_io_V_wire_en_0;
  wire[1:0] ArrayRowModule_2_io_H_out_22;
  wire[1:0] ArrayRowModule_2_io_H_out_21;
  wire[1:0] ArrayRowModule_2_io_H_out_20;
  wire[1:0] ArrayRowModule_2_io_H_out_19;
  wire[1:0] ArrayRowModule_2_io_H_out_18;
  wire[1:0] ArrayRowModule_2_io_H_out_17;
  wire[1:0] ArrayRowModule_2_io_H_out_16;
  wire[1:0] ArrayRowModule_2_io_H_out_15;
  wire[1:0] ArrayRowModule_2_io_H_out_14;
  wire[1:0] ArrayRowModule_2_io_H_out_13;
  wire[1:0] ArrayRowModule_2_io_H_out_12;
  wire[1:0] ArrayRowModule_2_io_H_out_11;
  wire[1:0] ArrayRowModule_2_io_H_out_10;
  wire[1:0] ArrayRowModule_2_io_H_out_9;
  wire[1:0] ArrayRowModule_2_io_H_out_8;
  wire[1:0] ArrayRowModule_2_io_H_out_7;
  wire[1:0] ArrayRowModule_2_io_H_out_6;
  wire[1:0] ArrayRowModule_2_io_H_out_5;
  wire[1:0] ArrayRowModule_2_io_H_out_4;
  wire[1:0] ArrayRowModule_2_io_H_out_3;
  wire[1:0] ArrayRowModule_2_io_H_out_2;
  wire[1:0] ArrayRowModule_2_io_H_out_1;
  wire[1:0] ArrayRowModule_2_io_H_out_0;
  wire[1:0] ArrayRowModule_2_io_G_wire_below_3;
  wire[1:0] ArrayRowModule_2_io_G_wire_below_2;
  wire[1:0] ArrayRowModule_2_io_G_wire_below_1;
  wire[1:0] ArrayRowModule_2_io_G_wire_below_0;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_32;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_31;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_30;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_29;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_28;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_27;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_26;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_25;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_24;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_23;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_22;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_21;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_20;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_19;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_18;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_17;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_16;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_15;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_14;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_13;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_12;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_11;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_10;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_9;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_8;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_7;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_6;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_5;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_4;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_3;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_2;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_1;
  wire[1:0] ArrayRowModule_2_io_H_wire_below_0;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_23;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_22;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_21;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_20;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_19;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_18;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_17;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_16;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_15;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_14;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_13;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_12;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_11;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_10;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_9;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_8;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_7;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_6;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_5;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_4;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_3;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_2;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_1;
  wire[1:0] ArrayRowModule_2_io_mem_bus_out_0;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_367;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_366;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_365;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_364;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_363;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_362;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_361;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_360;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_359;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_358;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_357;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_356;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_355;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_354;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_353;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_352;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_351;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_350;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_349;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_348;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_347;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_346;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_345;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_344;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_343;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_342;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_341;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_340;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_339;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_338;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_337;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_336;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_335;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_334;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_333;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_332;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_331;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_330;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_329;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_328;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_327;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_326;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_325;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_324;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_323;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_322;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_321;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_320;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_319;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_318;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_317;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_316;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_315;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_314;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_313;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_312;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_311;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_310;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_309;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_308;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_307;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_306;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_305;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_304;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_303;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_302;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_301;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_300;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_299;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_298;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_297;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_296;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_295;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_294;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_293;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_292;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_291;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_290;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_289;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_288;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_287;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_286;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_285;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_284;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_283;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_282;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_281;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_280;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_279;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_278;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_277;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_276;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_275;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_274;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_273;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_272;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_271;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_270;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_269;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_268;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_267;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_266;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_265;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_264;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_263;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_262;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_261;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_260;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_259;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_258;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_257;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_256;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_255;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_254;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_253;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_252;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_251;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_250;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_249;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_248;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_247;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_246;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_245;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_244;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_243;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_242;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_241;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_240;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_239;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_238;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_237;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_236;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_235;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_234;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_233;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_232;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_231;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_230;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_229;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_228;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_227;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_226;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_225;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_224;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_223;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_222;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_221;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_220;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_219;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_218;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_217;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_216;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_215;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_214;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_213;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_212;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_211;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_210;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_209;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_208;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_207;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_206;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_205;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_204;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_203;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_202;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_201;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_200;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_199;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_198;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_197;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_196;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_195;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_194;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_193;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_192;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_191;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_190;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_189;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_188;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_187;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_186;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_185;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_184;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_183;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_182;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_181;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_180;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_179;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_178;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_177;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_176;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_175;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_174;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_173;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_172;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_171;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_170;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_169;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_168;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_167;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_166;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_165;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_164;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_163;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_162;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_161;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_160;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_159;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_158;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_157;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_156;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_155;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_154;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_153;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_152;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_151;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_150;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_149;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_148;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_147;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_146;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_145;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_144;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_143;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_142;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_141;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_140;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_139;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_138;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_137;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_136;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_135;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_134;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_133;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_132;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_131;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_130;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_129;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_128;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_127;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_126;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_125;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_124;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_123;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_122;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_121;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_120;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_119;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_118;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_117;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_116;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_115;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_114;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_113;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_112;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_111;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_110;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_109;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_108;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_107;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_106;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_105;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_104;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_103;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_102;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_101;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_100;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_99;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_98;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_97;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_96;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_95;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_94;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_93;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_92;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_91;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_90;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_89;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_88;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_87;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_86;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_85;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_84;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_83;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_82;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_81;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_80;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_79;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_78;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_77;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_76;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_75;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_74;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_73;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_72;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_71;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_70;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_69;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_68;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_67;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_66;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_65;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_64;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_63;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_62;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_61;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_60;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_59;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_58;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_57;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_56;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_55;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_54;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_53;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_52;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_51;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_50;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_49;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_48;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_47;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_46;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_45;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_44;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_43;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_42;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_41;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_40;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_39;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_38;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_37;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_36;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_35;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_34;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_33;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_32;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_31;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_30;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_29;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_28;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_27;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_26;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_25;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_24;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_23;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_22;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_21;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_20;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_19;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_18;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_17;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_16;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_15;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_14;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_13;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_12;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_11;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_10;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_9;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_8;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_7;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_6;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_5;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_4;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_3;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_2;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_1;
  wire[1:0] ArrayRowModule_3_io_V_wire_out_0;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_22;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_21;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_20;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_19;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_18;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_17;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_16;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_15;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_14;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_13;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_12;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_11;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_10;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_9;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_8;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_7;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_6;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_5;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_4;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_3;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_2;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_1;
  wire[15:0] ArrayRowModule_3_io_V_wire_en_0;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_23;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_22;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_21;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_20;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_19;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_18;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_17;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_16;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_15;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_14;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_13;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_12;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_11;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_10;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_9;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_8;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_7;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_6;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_5;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_4;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_3;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_2;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_1;
  wire[1:0] ArrayRowModule_3_io_mem_bus_out_0;
  wire[1:0] VwireModule_io_VwirePorts_3_22_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_22_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_21_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_20_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_19_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_18_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_17_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_16_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_15_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_14_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_13_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_12_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_11_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_10_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_9_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_8_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_7_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_6_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_5_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_4_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_3_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_2_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_1_0_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_15_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_14_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_13_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_12_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_11_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_10_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_9_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_8_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_7_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_6_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_5_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_4_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_3_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_2_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_1_out;
  wire[1:0] VwireModule_io_VwirePorts_3_0_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_22_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_21_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_20_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_19_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_18_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_17_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_16_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_15_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_14_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_13_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_12_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_11_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_10_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_9_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_8_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_7_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_6_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_5_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_4_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_3_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_2_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_1_0_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_15_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_14_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_13_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_12_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_11_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_10_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_9_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_8_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_7_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_6_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_5_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_4_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_3_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_2_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_1_out;
  wire[1:0] VwireModule_io_VwirePorts_2_0_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_22_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_21_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_20_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_19_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_18_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_17_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_16_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_15_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_14_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_13_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_12_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_11_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_10_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_9_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_8_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_7_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_6_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_5_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_4_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_3_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_2_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_1_0_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_15_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_14_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_13_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_12_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_11_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_10_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_9_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_8_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_7_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_6_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_5_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_4_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_3_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_2_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_1_out;
  wire[1:0] VwireModule_io_VwirePorts_1_0_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_22_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_21_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_20_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_19_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_18_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_17_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_16_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_15_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_14_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_13_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_12_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_11_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_10_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_9_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_8_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_7_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_6_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_5_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_4_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_3_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_2_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_1_0_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_15_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_14_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_13_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_12_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_11_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_10_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_9_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_8_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_7_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_6_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_5_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_4_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_3_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_2_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_1_out;
  wire[1:0] VwireModule_io_VwirePorts_0_0_0_out;


`ifndef SYNTHESIS
// synthesis translate_off
  assign T1476 = {1{$random}};
  assign T1477 = {1{$random}};
  assign T1478 = {1{$random}};
  assign T1479 = {1{$random}};
  assign T1480 = {1{$random}};
  assign T1481 = {1{$random}};
  assign T1482 = {1{$random}};
  assign T1483 = {1{$random}};
  assign T1484 = {1{$random}};
  assign T1485 = {1{$random}};
  assign T1486 = {1{$random}};
  assign T1487 = {1{$random}};
  assign T1488 = {1{$random}};
  assign T1489 = {1{$random}};
  assign T1490 = {1{$random}};
  assign T1491 = {1{$random}};
  assign T1492 = {1{$random}};
  assign T1493 = {1{$random}};
  assign T1494 = {1{$random}};
  assign T1495 = {1{$random}};
  assign T1496 = {1{$random}};
  assign T1497 = {1{$random}};
  assign T1498 = {1{$random}};
  assign T1499 = {1{$random}};
  assign T1500 = {1{$random}};
  assign T1501 = {1{$random}};
  assign T1502 = {1{$random}};
  assign T1503 = {1{$random}};
  assign T1504 = {1{$random}};
  assign T1505 = {1{$random}};
  assign T1506 = {1{$random}};
  assign T1507 = {1{$random}};
  assign T1508 = {1{$random}};
  assign T1509 = {1{$random}};
  assign T1510 = {1{$random}};
  assign T1511 = {1{$random}};
  assign T1512 = {1{$random}};
  assign T1513 = {1{$random}};
  assign T1514 = {1{$random}};
  assign T1515 = {1{$random}};
  assign T1516 = {1{$random}};
  assign T1517 = {1{$random}};
  assign T1518 = {1{$random}};
  assign T1519 = {1{$random}};
  assign T1520 = {1{$random}};
  assign T1521 = {1{$random}};
  assign T1522 = {1{$random}};
  assign T1523 = {1{$random}};
  assign T1524 = {1{$random}};
  assign T1525 = {1{$random}};
  assign T1526 = {1{$random}};
  assign T1527 = {1{$random}};
  assign T1528 = {1{$random}};
  assign T1529 = {1{$random}};
  assign T1530 = {1{$random}};
  assign T1531 = {1{$random}};
  assign T1532 = {1{$random}};
  assign T1533 = {1{$random}};
  assign T1534 = {1{$random}};
  assign T1535 = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = ArrayRowModule_io_V_wire_en_0[1'h0];
  assign T1 = ArrayRowModule_io_V_wire_en_0[1'h1];
  assign T2 = ArrayRowModule_io_V_wire_en_0[2'h2];
  assign T3 = ArrayRowModule_io_V_wire_en_0[2'h3];
  assign T4 = ArrayRowModule_io_V_wire_en_0[3'h4];
  assign T5 = ArrayRowModule_io_V_wire_en_0[3'h5];
  assign T6 = ArrayRowModule_io_V_wire_en_0[3'h6];
  assign T7 = ArrayRowModule_io_V_wire_en_0[3'h7];
  assign T8 = ArrayRowModule_io_V_wire_en_0[4'h8];
  assign T9 = ArrayRowModule_io_V_wire_en_0[4'h9];
  assign T10 = ArrayRowModule_io_V_wire_en_0[4'ha];
  assign T11 = ArrayRowModule_io_V_wire_en_0[4'hb];
  assign T12 = ArrayRowModule_io_V_wire_en_0[4'hc];
  assign T13 = ArrayRowModule_io_V_wire_en_0[4'hd];
  assign T14 = ArrayRowModule_io_V_wire_en_0[4'he];
  assign T15 = ArrayRowModule_io_V_wire_en_0[4'hf];
  assign T16 = ArrayRowModule_io_V_wire_en_1[1'h0];
  assign T17 = ArrayRowModule_io_V_wire_en_1[1'h1];
  assign T18 = ArrayRowModule_io_V_wire_en_1[2'h2];
  assign T19 = ArrayRowModule_io_V_wire_en_1[2'h3];
  assign T20 = ArrayRowModule_io_V_wire_en_1[3'h4];
  assign T21 = ArrayRowModule_io_V_wire_en_1[3'h5];
  assign T22 = ArrayRowModule_io_V_wire_en_1[3'h6];
  assign T23 = ArrayRowModule_io_V_wire_en_1[3'h7];
  assign T24 = ArrayRowModule_io_V_wire_en_1[4'h8];
  assign T25 = ArrayRowModule_io_V_wire_en_1[4'h9];
  assign T26 = ArrayRowModule_io_V_wire_en_1[4'ha];
  assign T27 = ArrayRowModule_io_V_wire_en_1[4'hb];
  assign T28 = ArrayRowModule_io_V_wire_en_1[4'hc];
  assign T29 = ArrayRowModule_io_V_wire_en_1[4'hd];
  assign T30 = ArrayRowModule_io_V_wire_en_1[4'he];
  assign T31 = ArrayRowModule_io_V_wire_en_1[4'hf];
  assign T32 = ArrayRowModule_io_V_wire_en_2[1'h0];
  assign T33 = ArrayRowModule_io_V_wire_en_2[1'h1];
  assign T34 = ArrayRowModule_io_V_wire_en_2[2'h2];
  assign T35 = ArrayRowModule_io_V_wire_en_2[2'h3];
  assign T36 = ArrayRowModule_io_V_wire_en_2[3'h4];
  assign T37 = ArrayRowModule_io_V_wire_en_2[3'h5];
  assign T38 = ArrayRowModule_io_V_wire_en_2[3'h6];
  assign T39 = ArrayRowModule_io_V_wire_en_2[3'h7];
  assign T40 = ArrayRowModule_io_V_wire_en_2[4'h8];
  assign T41 = ArrayRowModule_io_V_wire_en_2[4'h9];
  assign T42 = ArrayRowModule_io_V_wire_en_2[4'ha];
  assign T43 = ArrayRowModule_io_V_wire_en_2[4'hb];
  assign T44 = ArrayRowModule_io_V_wire_en_2[4'hc];
  assign T45 = ArrayRowModule_io_V_wire_en_2[4'hd];
  assign T46 = ArrayRowModule_io_V_wire_en_2[4'he];
  assign T47 = ArrayRowModule_io_V_wire_en_2[4'hf];
  assign T48 = ArrayRowModule_io_V_wire_en_3[1'h0];
  assign T49 = ArrayRowModule_io_V_wire_en_3[1'h1];
  assign T50 = ArrayRowModule_io_V_wire_en_3[2'h2];
  assign T51 = ArrayRowModule_io_V_wire_en_3[2'h3];
  assign T52 = ArrayRowModule_io_V_wire_en_3[3'h4];
  assign T53 = ArrayRowModule_io_V_wire_en_3[3'h5];
  assign T54 = ArrayRowModule_io_V_wire_en_3[3'h6];
  assign T55 = ArrayRowModule_io_V_wire_en_3[3'h7];
  assign T56 = ArrayRowModule_io_V_wire_en_3[4'h8];
  assign T57 = ArrayRowModule_io_V_wire_en_3[4'h9];
  assign T58 = ArrayRowModule_io_V_wire_en_3[4'ha];
  assign T59 = ArrayRowModule_io_V_wire_en_3[4'hb];
  assign T60 = ArrayRowModule_io_V_wire_en_3[4'hc];
  assign T61 = ArrayRowModule_io_V_wire_en_3[4'hd];
  assign T62 = ArrayRowModule_io_V_wire_en_3[4'he];
  assign T63 = ArrayRowModule_io_V_wire_en_3[4'hf];
  assign T64 = ArrayRowModule_io_V_wire_en_4[1'h0];
  assign T65 = ArrayRowModule_io_V_wire_en_4[1'h1];
  assign T66 = ArrayRowModule_io_V_wire_en_4[2'h2];
  assign T67 = ArrayRowModule_io_V_wire_en_4[2'h3];
  assign T68 = ArrayRowModule_io_V_wire_en_4[3'h4];
  assign T69 = ArrayRowModule_io_V_wire_en_4[3'h5];
  assign T70 = ArrayRowModule_io_V_wire_en_4[3'h6];
  assign T71 = ArrayRowModule_io_V_wire_en_4[3'h7];
  assign T72 = ArrayRowModule_io_V_wire_en_4[4'h8];
  assign T73 = ArrayRowModule_io_V_wire_en_4[4'h9];
  assign T74 = ArrayRowModule_io_V_wire_en_4[4'ha];
  assign T75 = ArrayRowModule_io_V_wire_en_4[4'hb];
  assign T76 = ArrayRowModule_io_V_wire_en_4[4'hc];
  assign T77 = ArrayRowModule_io_V_wire_en_4[4'hd];
  assign T78 = ArrayRowModule_io_V_wire_en_4[4'he];
  assign T79 = ArrayRowModule_io_V_wire_en_4[4'hf];
  assign T80 = ArrayRowModule_io_V_wire_en_5[1'h0];
  assign T81 = ArrayRowModule_io_V_wire_en_5[1'h1];
  assign T82 = ArrayRowModule_io_V_wire_en_5[2'h2];
  assign T83 = ArrayRowModule_io_V_wire_en_5[2'h3];
  assign T84 = ArrayRowModule_io_V_wire_en_5[3'h4];
  assign T85 = ArrayRowModule_io_V_wire_en_5[3'h5];
  assign T86 = ArrayRowModule_io_V_wire_en_5[3'h6];
  assign T87 = ArrayRowModule_io_V_wire_en_5[3'h7];
  assign T88 = ArrayRowModule_io_V_wire_en_5[4'h8];
  assign T89 = ArrayRowModule_io_V_wire_en_5[4'h9];
  assign T90 = ArrayRowModule_io_V_wire_en_5[4'ha];
  assign T91 = ArrayRowModule_io_V_wire_en_5[4'hb];
  assign T92 = ArrayRowModule_io_V_wire_en_5[4'hc];
  assign T93 = ArrayRowModule_io_V_wire_en_5[4'hd];
  assign T94 = ArrayRowModule_io_V_wire_en_5[4'he];
  assign T95 = ArrayRowModule_io_V_wire_en_5[4'hf];
  assign T96 = ArrayRowModule_io_V_wire_en_6[1'h0];
  assign T97 = ArrayRowModule_io_V_wire_en_6[1'h1];
  assign T98 = ArrayRowModule_io_V_wire_en_6[2'h2];
  assign T99 = ArrayRowModule_io_V_wire_en_6[2'h3];
  assign T100 = ArrayRowModule_io_V_wire_en_6[3'h4];
  assign T101 = ArrayRowModule_io_V_wire_en_6[3'h5];
  assign T102 = ArrayRowModule_io_V_wire_en_6[3'h6];
  assign T103 = ArrayRowModule_io_V_wire_en_6[3'h7];
  assign T104 = ArrayRowModule_io_V_wire_en_6[4'h8];
  assign T105 = ArrayRowModule_io_V_wire_en_6[4'h9];
  assign T106 = ArrayRowModule_io_V_wire_en_6[4'ha];
  assign T107 = ArrayRowModule_io_V_wire_en_6[4'hb];
  assign T108 = ArrayRowModule_io_V_wire_en_6[4'hc];
  assign T109 = ArrayRowModule_io_V_wire_en_6[4'hd];
  assign T110 = ArrayRowModule_io_V_wire_en_6[4'he];
  assign T111 = ArrayRowModule_io_V_wire_en_6[4'hf];
  assign T112 = ArrayRowModule_io_V_wire_en_7[1'h0];
  assign T113 = ArrayRowModule_io_V_wire_en_7[1'h1];
  assign T114 = ArrayRowModule_io_V_wire_en_7[2'h2];
  assign T115 = ArrayRowModule_io_V_wire_en_7[2'h3];
  assign T116 = ArrayRowModule_io_V_wire_en_7[3'h4];
  assign T117 = ArrayRowModule_io_V_wire_en_7[3'h5];
  assign T118 = ArrayRowModule_io_V_wire_en_7[3'h6];
  assign T119 = ArrayRowModule_io_V_wire_en_7[3'h7];
  assign T120 = ArrayRowModule_io_V_wire_en_7[4'h8];
  assign T121 = ArrayRowModule_io_V_wire_en_7[4'h9];
  assign T122 = ArrayRowModule_io_V_wire_en_7[4'ha];
  assign T123 = ArrayRowModule_io_V_wire_en_7[4'hb];
  assign T124 = ArrayRowModule_io_V_wire_en_7[4'hc];
  assign T125 = ArrayRowModule_io_V_wire_en_7[4'hd];
  assign T126 = ArrayRowModule_io_V_wire_en_7[4'he];
  assign T127 = ArrayRowModule_io_V_wire_en_7[4'hf];
  assign T128 = ArrayRowModule_io_V_wire_en_8[1'h0];
  assign T129 = ArrayRowModule_io_V_wire_en_8[1'h1];
  assign T130 = ArrayRowModule_io_V_wire_en_8[2'h2];
  assign T131 = ArrayRowModule_io_V_wire_en_8[2'h3];
  assign T132 = ArrayRowModule_io_V_wire_en_8[3'h4];
  assign T133 = ArrayRowModule_io_V_wire_en_8[3'h5];
  assign T134 = ArrayRowModule_io_V_wire_en_8[3'h6];
  assign T135 = ArrayRowModule_io_V_wire_en_8[3'h7];
  assign T136 = ArrayRowModule_io_V_wire_en_8[4'h8];
  assign T137 = ArrayRowModule_io_V_wire_en_8[4'h9];
  assign T138 = ArrayRowModule_io_V_wire_en_8[4'ha];
  assign T139 = ArrayRowModule_io_V_wire_en_8[4'hb];
  assign T140 = ArrayRowModule_io_V_wire_en_8[4'hc];
  assign T141 = ArrayRowModule_io_V_wire_en_8[4'hd];
  assign T142 = ArrayRowModule_io_V_wire_en_8[4'he];
  assign T143 = ArrayRowModule_io_V_wire_en_8[4'hf];
  assign T144 = ArrayRowModule_io_V_wire_en_9[1'h0];
  assign T145 = ArrayRowModule_io_V_wire_en_9[1'h1];
  assign T146 = ArrayRowModule_io_V_wire_en_9[2'h2];
  assign T147 = ArrayRowModule_io_V_wire_en_9[2'h3];
  assign T148 = ArrayRowModule_io_V_wire_en_9[3'h4];
  assign T149 = ArrayRowModule_io_V_wire_en_9[3'h5];
  assign T150 = ArrayRowModule_io_V_wire_en_9[3'h6];
  assign T151 = ArrayRowModule_io_V_wire_en_9[3'h7];
  assign T152 = ArrayRowModule_io_V_wire_en_9[4'h8];
  assign T153 = ArrayRowModule_io_V_wire_en_9[4'h9];
  assign T154 = ArrayRowModule_io_V_wire_en_9[4'ha];
  assign T155 = ArrayRowModule_io_V_wire_en_9[4'hb];
  assign T156 = ArrayRowModule_io_V_wire_en_9[4'hc];
  assign T157 = ArrayRowModule_io_V_wire_en_9[4'hd];
  assign T158 = ArrayRowModule_io_V_wire_en_9[4'he];
  assign T159 = ArrayRowModule_io_V_wire_en_9[4'hf];
  assign T160 = ArrayRowModule_io_V_wire_en_10[1'h0];
  assign T161 = ArrayRowModule_io_V_wire_en_10[1'h1];
  assign T162 = ArrayRowModule_io_V_wire_en_10[2'h2];
  assign T163 = ArrayRowModule_io_V_wire_en_10[2'h3];
  assign T164 = ArrayRowModule_io_V_wire_en_10[3'h4];
  assign T165 = ArrayRowModule_io_V_wire_en_10[3'h5];
  assign T166 = ArrayRowModule_io_V_wire_en_10[3'h6];
  assign T167 = ArrayRowModule_io_V_wire_en_10[3'h7];
  assign T168 = ArrayRowModule_io_V_wire_en_10[4'h8];
  assign T169 = ArrayRowModule_io_V_wire_en_10[4'h9];
  assign T170 = ArrayRowModule_io_V_wire_en_10[4'ha];
  assign T171 = ArrayRowModule_io_V_wire_en_10[4'hb];
  assign T172 = ArrayRowModule_io_V_wire_en_10[4'hc];
  assign T173 = ArrayRowModule_io_V_wire_en_10[4'hd];
  assign T174 = ArrayRowModule_io_V_wire_en_10[4'he];
  assign T175 = ArrayRowModule_io_V_wire_en_10[4'hf];
  assign T176 = ArrayRowModule_io_V_wire_en_11[1'h0];
  assign T177 = ArrayRowModule_io_V_wire_en_11[1'h1];
  assign T178 = ArrayRowModule_io_V_wire_en_11[2'h2];
  assign T179 = ArrayRowModule_io_V_wire_en_11[2'h3];
  assign T180 = ArrayRowModule_io_V_wire_en_11[3'h4];
  assign T181 = ArrayRowModule_io_V_wire_en_11[3'h5];
  assign T182 = ArrayRowModule_io_V_wire_en_11[3'h6];
  assign T183 = ArrayRowModule_io_V_wire_en_11[3'h7];
  assign T184 = ArrayRowModule_io_V_wire_en_11[4'h8];
  assign T185 = ArrayRowModule_io_V_wire_en_11[4'h9];
  assign T186 = ArrayRowModule_io_V_wire_en_11[4'ha];
  assign T187 = ArrayRowModule_io_V_wire_en_11[4'hb];
  assign T188 = ArrayRowModule_io_V_wire_en_11[4'hc];
  assign T189 = ArrayRowModule_io_V_wire_en_11[4'hd];
  assign T190 = ArrayRowModule_io_V_wire_en_11[4'he];
  assign T191 = ArrayRowModule_io_V_wire_en_11[4'hf];
  assign T192 = ArrayRowModule_io_V_wire_en_12[1'h0];
  assign T193 = ArrayRowModule_io_V_wire_en_12[1'h1];
  assign T194 = ArrayRowModule_io_V_wire_en_12[2'h2];
  assign T195 = ArrayRowModule_io_V_wire_en_12[2'h3];
  assign T196 = ArrayRowModule_io_V_wire_en_12[3'h4];
  assign T197 = ArrayRowModule_io_V_wire_en_12[3'h5];
  assign T198 = ArrayRowModule_io_V_wire_en_12[3'h6];
  assign T199 = ArrayRowModule_io_V_wire_en_12[3'h7];
  assign T200 = ArrayRowModule_io_V_wire_en_12[4'h8];
  assign T201 = ArrayRowModule_io_V_wire_en_12[4'h9];
  assign T202 = ArrayRowModule_io_V_wire_en_12[4'ha];
  assign T203 = ArrayRowModule_io_V_wire_en_12[4'hb];
  assign T204 = ArrayRowModule_io_V_wire_en_12[4'hc];
  assign T205 = ArrayRowModule_io_V_wire_en_12[4'hd];
  assign T206 = ArrayRowModule_io_V_wire_en_12[4'he];
  assign T207 = ArrayRowModule_io_V_wire_en_12[4'hf];
  assign T208 = ArrayRowModule_io_V_wire_en_13[1'h0];
  assign T209 = ArrayRowModule_io_V_wire_en_13[1'h1];
  assign T210 = ArrayRowModule_io_V_wire_en_13[2'h2];
  assign T211 = ArrayRowModule_io_V_wire_en_13[2'h3];
  assign T212 = ArrayRowModule_io_V_wire_en_13[3'h4];
  assign T213 = ArrayRowModule_io_V_wire_en_13[3'h5];
  assign T214 = ArrayRowModule_io_V_wire_en_13[3'h6];
  assign T215 = ArrayRowModule_io_V_wire_en_13[3'h7];
  assign T216 = ArrayRowModule_io_V_wire_en_13[4'h8];
  assign T217 = ArrayRowModule_io_V_wire_en_13[4'h9];
  assign T218 = ArrayRowModule_io_V_wire_en_13[4'ha];
  assign T219 = ArrayRowModule_io_V_wire_en_13[4'hb];
  assign T220 = ArrayRowModule_io_V_wire_en_13[4'hc];
  assign T221 = ArrayRowModule_io_V_wire_en_13[4'hd];
  assign T222 = ArrayRowModule_io_V_wire_en_13[4'he];
  assign T223 = ArrayRowModule_io_V_wire_en_13[4'hf];
  assign T224 = ArrayRowModule_io_V_wire_en_14[1'h0];
  assign T225 = ArrayRowModule_io_V_wire_en_14[1'h1];
  assign T226 = ArrayRowModule_io_V_wire_en_14[2'h2];
  assign T227 = ArrayRowModule_io_V_wire_en_14[2'h3];
  assign T228 = ArrayRowModule_io_V_wire_en_14[3'h4];
  assign T229 = ArrayRowModule_io_V_wire_en_14[3'h5];
  assign T230 = ArrayRowModule_io_V_wire_en_14[3'h6];
  assign T231 = ArrayRowModule_io_V_wire_en_14[3'h7];
  assign T232 = ArrayRowModule_io_V_wire_en_14[4'h8];
  assign T233 = ArrayRowModule_io_V_wire_en_14[4'h9];
  assign T234 = ArrayRowModule_io_V_wire_en_14[4'ha];
  assign T235 = ArrayRowModule_io_V_wire_en_14[4'hb];
  assign T236 = ArrayRowModule_io_V_wire_en_14[4'hc];
  assign T237 = ArrayRowModule_io_V_wire_en_14[4'hd];
  assign T238 = ArrayRowModule_io_V_wire_en_14[4'he];
  assign T239 = ArrayRowModule_io_V_wire_en_14[4'hf];
  assign T240 = ArrayRowModule_io_V_wire_en_15[1'h0];
  assign T241 = ArrayRowModule_io_V_wire_en_15[1'h1];
  assign T242 = ArrayRowModule_io_V_wire_en_15[2'h2];
  assign T243 = ArrayRowModule_io_V_wire_en_15[2'h3];
  assign T244 = ArrayRowModule_io_V_wire_en_15[3'h4];
  assign T245 = ArrayRowModule_io_V_wire_en_15[3'h5];
  assign T246 = ArrayRowModule_io_V_wire_en_15[3'h6];
  assign T247 = ArrayRowModule_io_V_wire_en_15[3'h7];
  assign T248 = ArrayRowModule_io_V_wire_en_15[4'h8];
  assign T249 = ArrayRowModule_io_V_wire_en_15[4'h9];
  assign T250 = ArrayRowModule_io_V_wire_en_15[4'ha];
  assign T251 = ArrayRowModule_io_V_wire_en_15[4'hb];
  assign T252 = ArrayRowModule_io_V_wire_en_15[4'hc];
  assign T253 = ArrayRowModule_io_V_wire_en_15[4'hd];
  assign T254 = ArrayRowModule_io_V_wire_en_15[4'he];
  assign T255 = ArrayRowModule_io_V_wire_en_15[4'hf];
  assign T256 = ArrayRowModule_io_V_wire_en_16[1'h0];
  assign T257 = ArrayRowModule_io_V_wire_en_16[1'h1];
  assign T258 = ArrayRowModule_io_V_wire_en_16[2'h2];
  assign T259 = ArrayRowModule_io_V_wire_en_16[2'h3];
  assign T260 = ArrayRowModule_io_V_wire_en_16[3'h4];
  assign T261 = ArrayRowModule_io_V_wire_en_16[3'h5];
  assign T262 = ArrayRowModule_io_V_wire_en_16[3'h6];
  assign T263 = ArrayRowModule_io_V_wire_en_16[3'h7];
  assign T264 = ArrayRowModule_io_V_wire_en_16[4'h8];
  assign T265 = ArrayRowModule_io_V_wire_en_16[4'h9];
  assign T266 = ArrayRowModule_io_V_wire_en_16[4'ha];
  assign T267 = ArrayRowModule_io_V_wire_en_16[4'hb];
  assign T268 = ArrayRowModule_io_V_wire_en_16[4'hc];
  assign T269 = ArrayRowModule_io_V_wire_en_16[4'hd];
  assign T270 = ArrayRowModule_io_V_wire_en_16[4'he];
  assign T271 = ArrayRowModule_io_V_wire_en_16[4'hf];
  assign T272 = ArrayRowModule_io_V_wire_en_17[1'h0];
  assign T273 = ArrayRowModule_io_V_wire_en_17[1'h1];
  assign T274 = ArrayRowModule_io_V_wire_en_17[2'h2];
  assign T275 = ArrayRowModule_io_V_wire_en_17[2'h3];
  assign T276 = ArrayRowModule_io_V_wire_en_17[3'h4];
  assign T277 = ArrayRowModule_io_V_wire_en_17[3'h5];
  assign T278 = ArrayRowModule_io_V_wire_en_17[3'h6];
  assign T279 = ArrayRowModule_io_V_wire_en_17[3'h7];
  assign T280 = ArrayRowModule_io_V_wire_en_17[4'h8];
  assign T281 = ArrayRowModule_io_V_wire_en_17[4'h9];
  assign T282 = ArrayRowModule_io_V_wire_en_17[4'ha];
  assign T283 = ArrayRowModule_io_V_wire_en_17[4'hb];
  assign T284 = ArrayRowModule_io_V_wire_en_17[4'hc];
  assign T285 = ArrayRowModule_io_V_wire_en_17[4'hd];
  assign T286 = ArrayRowModule_io_V_wire_en_17[4'he];
  assign T287 = ArrayRowModule_io_V_wire_en_17[4'hf];
  assign T288 = ArrayRowModule_io_V_wire_en_18[1'h0];
  assign T289 = ArrayRowModule_io_V_wire_en_18[1'h1];
  assign T290 = ArrayRowModule_io_V_wire_en_18[2'h2];
  assign T291 = ArrayRowModule_io_V_wire_en_18[2'h3];
  assign T292 = ArrayRowModule_io_V_wire_en_18[3'h4];
  assign T293 = ArrayRowModule_io_V_wire_en_18[3'h5];
  assign T294 = ArrayRowModule_io_V_wire_en_18[3'h6];
  assign T295 = ArrayRowModule_io_V_wire_en_18[3'h7];
  assign T296 = ArrayRowModule_io_V_wire_en_18[4'h8];
  assign T297 = ArrayRowModule_io_V_wire_en_18[4'h9];
  assign T298 = ArrayRowModule_io_V_wire_en_18[4'ha];
  assign T299 = ArrayRowModule_io_V_wire_en_18[4'hb];
  assign T300 = ArrayRowModule_io_V_wire_en_18[4'hc];
  assign T301 = ArrayRowModule_io_V_wire_en_18[4'hd];
  assign T302 = ArrayRowModule_io_V_wire_en_18[4'he];
  assign T303 = ArrayRowModule_io_V_wire_en_18[4'hf];
  assign T304 = ArrayRowModule_io_V_wire_en_19[1'h0];
  assign T305 = ArrayRowModule_io_V_wire_en_19[1'h1];
  assign T306 = ArrayRowModule_io_V_wire_en_19[2'h2];
  assign T307 = ArrayRowModule_io_V_wire_en_19[2'h3];
  assign T308 = ArrayRowModule_io_V_wire_en_19[3'h4];
  assign T309 = ArrayRowModule_io_V_wire_en_19[3'h5];
  assign T310 = ArrayRowModule_io_V_wire_en_19[3'h6];
  assign T311 = ArrayRowModule_io_V_wire_en_19[3'h7];
  assign T312 = ArrayRowModule_io_V_wire_en_19[4'h8];
  assign T313 = ArrayRowModule_io_V_wire_en_19[4'h9];
  assign T314 = ArrayRowModule_io_V_wire_en_19[4'ha];
  assign T315 = ArrayRowModule_io_V_wire_en_19[4'hb];
  assign T316 = ArrayRowModule_io_V_wire_en_19[4'hc];
  assign T317 = ArrayRowModule_io_V_wire_en_19[4'hd];
  assign T318 = ArrayRowModule_io_V_wire_en_19[4'he];
  assign T319 = ArrayRowModule_io_V_wire_en_19[4'hf];
  assign T320 = ArrayRowModule_io_V_wire_en_20[1'h0];
  assign T321 = ArrayRowModule_io_V_wire_en_20[1'h1];
  assign T322 = ArrayRowModule_io_V_wire_en_20[2'h2];
  assign T323 = ArrayRowModule_io_V_wire_en_20[2'h3];
  assign T324 = ArrayRowModule_io_V_wire_en_20[3'h4];
  assign T325 = ArrayRowModule_io_V_wire_en_20[3'h5];
  assign T326 = ArrayRowModule_io_V_wire_en_20[3'h6];
  assign T327 = ArrayRowModule_io_V_wire_en_20[3'h7];
  assign T328 = ArrayRowModule_io_V_wire_en_20[4'h8];
  assign T329 = ArrayRowModule_io_V_wire_en_20[4'h9];
  assign T330 = ArrayRowModule_io_V_wire_en_20[4'ha];
  assign T331 = ArrayRowModule_io_V_wire_en_20[4'hb];
  assign T332 = ArrayRowModule_io_V_wire_en_20[4'hc];
  assign T333 = ArrayRowModule_io_V_wire_en_20[4'hd];
  assign T334 = ArrayRowModule_io_V_wire_en_20[4'he];
  assign T335 = ArrayRowModule_io_V_wire_en_20[4'hf];
  assign T336 = ArrayRowModule_io_V_wire_en_21[1'h0];
  assign T337 = ArrayRowModule_io_V_wire_en_21[1'h1];
  assign T338 = ArrayRowModule_io_V_wire_en_21[2'h2];
  assign T339 = ArrayRowModule_io_V_wire_en_21[2'h3];
  assign T340 = ArrayRowModule_io_V_wire_en_21[3'h4];
  assign T341 = ArrayRowModule_io_V_wire_en_21[3'h5];
  assign T342 = ArrayRowModule_io_V_wire_en_21[3'h6];
  assign T343 = ArrayRowModule_io_V_wire_en_21[3'h7];
  assign T344 = ArrayRowModule_io_V_wire_en_21[4'h8];
  assign T345 = ArrayRowModule_io_V_wire_en_21[4'h9];
  assign T346 = ArrayRowModule_io_V_wire_en_21[4'ha];
  assign T347 = ArrayRowModule_io_V_wire_en_21[4'hb];
  assign T348 = ArrayRowModule_io_V_wire_en_21[4'hc];
  assign T349 = ArrayRowModule_io_V_wire_en_21[4'hd];
  assign T350 = ArrayRowModule_io_V_wire_en_21[4'he];
  assign T351 = ArrayRowModule_io_V_wire_en_21[4'hf];
  assign T352 = ArrayRowModule_io_V_wire_en_22[1'h0];
  assign T353 = ArrayRowModule_io_V_wire_en_22[1'h1];
  assign T354 = ArrayRowModule_io_V_wire_en_22[2'h2];
  assign T355 = ArrayRowModule_io_V_wire_en_22[2'h3];
  assign T356 = ArrayRowModule_io_V_wire_en_22[3'h4];
  assign T357 = ArrayRowModule_io_V_wire_en_22[3'h5];
  assign T358 = ArrayRowModule_io_V_wire_en_22[3'h6];
  assign T359 = ArrayRowModule_io_V_wire_en_22[3'h7];
  assign T360 = ArrayRowModule_io_V_wire_en_22[4'h8];
  assign T361 = ArrayRowModule_io_V_wire_en_22[4'h9];
  assign T362 = ArrayRowModule_io_V_wire_en_22[4'ha];
  assign T363 = ArrayRowModule_io_V_wire_en_22[4'hb];
  assign T364 = ArrayRowModule_io_V_wire_en_22[4'hc];
  assign T365 = ArrayRowModule_io_V_wire_en_22[4'hd];
  assign T366 = ArrayRowModule_io_V_wire_en_22[4'he];
  assign T367 = ArrayRowModule_io_V_wire_en_22[4'hf];
  assign T368 = ArrayRowModule_1_io_V_wire_en_0[1'h0];
  assign T369 = ArrayRowModule_1_io_V_wire_en_0[1'h1];
  assign T370 = ArrayRowModule_1_io_V_wire_en_0[2'h2];
  assign T371 = ArrayRowModule_1_io_V_wire_en_0[2'h3];
  assign T372 = ArrayRowModule_1_io_V_wire_en_0[3'h4];
  assign T373 = ArrayRowModule_1_io_V_wire_en_0[3'h5];
  assign T374 = ArrayRowModule_1_io_V_wire_en_0[3'h6];
  assign T375 = ArrayRowModule_1_io_V_wire_en_0[3'h7];
  assign T376 = ArrayRowModule_1_io_V_wire_en_0[4'h8];
  assign T377 = ArrayRowModule_1_io_V_wire_en_0[4'h9];
  assign T378 = ArrayRowModule_1_io_V_wire_en_0[4'ha];
  assign T379 = ArrayRowModule_1_io_V_wire_en_0[4'hb];
  assign T380 = ArrayRowModule_1_io_V_wire_en_0[4'hc];
  assign T381 = ArrayRowModule_1_io_V_wire_en_0[4'hd];
  assign T382 = ArrayRowModule_1_io_V_wire_en_0[4'he];
  assign T383 = ArrayRowModule_1_io_V_wire_en_0[4'hf];
  assign T384 = ArrayRowModule_1_io_V_wire_en_1[1'h0];
  assign T385 = ArrayRowModule_1_io_V_wire_en_1[1'h1];
  assign T386 = ArrayRowModule_1_io_V_wire_en_1[2'h2];
  assign T387 = ArrayRowModule_1_io_V_wire_en_1[2'h3];
  assign T388 = ArrayRowModule_1_io_V_wire_en_1[3'h4];
  assign T389 = ArrayRowModule_1_io_V_wire_en_1[3'h5];
  assign T390 = ArrayRowModule_1_io_V_wire_en_1[3'h6];
  assign T391 = ArrayRowModule_1_io_V_wire_en_1[3'h7];
  assign T392 = ArrayRowModule_1_io_V_wire_en_1[4'h8];
  assign T393 = ArrayRowModule_1_io_V_wire_en_1[4'h9];
  assign T394 = ArrayRowModule_1_io_V_wire_en_1[4'ha];
  assign T395 = ArrayRowModule_1_io_V_wire_en_1[4'hb];
  assign T396 = ArrayRowModule_1_io_V_wire_en_1[4'hc];
  assign T397 = ArrayRowModule_1_io_V_wire_en_1[4'hd];
  assign T398 = ArrayRowModule_1_io_V_wire_en_1[4'he];
  assign T399 = ArrayRowModule_1_io_V_wire_en_1[4'hf];
  assign T400 = ArrayRowModule_1_io_V_wire_en_2[1'h0];
  assign T401 = ArrayRowModule_1_io_V_wire_en_2[1'h1];
  assign T402 = ArrayRowModule_1_io_V_wire_en_2[2'h2];
  assign T403 = ArrayRowModule_1_io_V_wire_en_2[2'h3];
  assign T404 = ArrayRowModule_1_io_V_wire_en_2[3'h4];
  assign T405 = ArrayRowModule_1_io_V_wire_en_2[3'h5];
  assign T406 = ArrayRowModule_1_io_V_wire_en_2[3'h6];
  assign T407 = ArrayRowModule_1_io_V_wire_en_2[3'h7];
  assign T408 = ArrayRowModule_1_io_V_wire_en_2[4'h8];
  assign T409 = ArrayRowModule_1_io_V_wire_en_2[4'h9];
  assign T410 = ArrayRowModule_1_io_V_wire_en_2[4'ha];
  assign T411 = ArrayRowModule_1_io_V_wire_en_2[4'hb];
  assign T412 = ArrayRowModule_1_io_V_wire_en_2[4'hc];
  assign T413 = ArrayRowModule_1_io_V_wire_en_2[4'hd];
  assign T414 = ArrayRowModule_1_io_V_wire_en_2[4'he];
  assign T415 = ArrayRowModule_1_io_V_wire_en_2[4'hf];
  assign T416 = ArrayRowModule_1_io_V_wire_en_3[1'h0];
  assign T417 = ArrayRowModule_1_io_V_wire_en_3[1'h1];
  assign T418 = ArrayRowModule_1_io_V_wire_en_3[2'h2];
  assign T419 = ArrayRowModule_1_io_V_wire_en_3[2'h3];
  assign T420 = ArrayRowModule_1_io_V_wire_en_3[3'h4];
  assign T421 = ArrayRowModule_1_io_V_wire_en_3[3'h5];
  assign T422 = ArrayRowModule_1_io_V_wire_en_3[3'h6];
  assign T423 = ArrayRowModule_1_io_V_wire_en_3[3'h7];
  assign T424 = ArrayRowModule_1_io_V_wire_en_3[4'h8];
  assign T425 = ArrayRowModule_1_io_V_wire_en_3[4'h9];
  assign T426 = ArrayRowModule_1_io_V_wire_en_3[4'ha];
  assign T427 = ArrayRowModule_1_io_V_wire_en_3[4'hb];
  assign T428 = ArrayRowModule_1_io_V_wire_en_3[4'hc];
  assign T429 = ArrayRowModule_1_io_V_wire_en_3[4'hd];
  assign T430 = ArrayRowModule_1_io_V_wire_en_3[4'he];
  assign T431 = ArrayRowModule_1_io_V_wire_en_3[4'hf];
  assign T432 = ArrayRowModule_1_io_V_wire_en_4[1'h0];
  assign T433 = ArrayRowModule_1_io_V_wire_en_4[1'h1];
  assign T434 = ArrayRowModule_1_io_V_wire_en_4[2'h2];
  assign T435 = ArrayRowModule_1_io_V_wire_en_4[2'h3];
  assign T436 = ArrayRowModule_1_io_V_wire_en_4[3'h4];
  assign T437 = ArrayRowModule_1_io_V_wire_en_4[3'h5];
  assign T438 = ArrayRowModule_1_io_V_wire_en_4[3'h6];
  assign T439 = ArrayRowModule_1_io_V_wire_en_4[3'h7];
  assign T440 = ArrayRowModule_1_io_V_wire_en_4[4'h8];
  assign T441 = ArrayRowModule_1_io_V_wire_en_4[4'h9];
  assign T442 = ArrayRowModule_1_io_V_wire_en_4[4'ha];
  assign T443 = ArrayRowModule_1_io_V_wire_en_4[4'hb];
  assign T444 = ArrayRowModule_1_io_V_wire_en_4[4'hc];
  assign T445 = ArrayRowModule_1_io_V_wire_en_4[4'hd];
  assign T446 = ArrayRowModule_1_io_V_wire_en_4[4'he];
  assign T447 = ArrayRowModule_1_io_V_wire_en_4[4'hf];
  assign T448 = ArrayRowModule_1_io_V_wire_en_5[1'h0];
  assign T449 = ArrayRowModule_1_io_V_wire_en_5[1'h1];
  assign T450 = ArrayRowModule_1_io_V_wire_en_5[2'h2];
  assign T451 = ArrayRowModule_1_io_V_wire_en_5[2'h3];
  assign T452 = ArrayRowModule_1_io_V_wire_en_5[3'h4];
  assign T453 = ArrayRowModule_1_io_V_wire_en_5[3'h5];
  assign T454 = ArrayRowModule_1_io_V_wire_en_5[3'h6];
  assign T455 = ArrayRowModule_1_io_V_wire_en_5[3'h7];
  assign T456 = ArrayRowModule_1_io_V_wire_en_5[4'h8];
  assign T457 = ArrayRowModule_1_io_V_wire_en_5[4'h9];
  assign T458 = ArrayRowModule_1_io_V_wire_en_5[4'ha];
  assign T459 = ArrayRowModule_1_io_V_wire_en_5[4'hb];
  assign T460 = ArrayRowModule_1_io_V_wire_en_5[4'hc];
  assign T461 = ArrayRowModule_1_io_V_wire_en_5[4'hd];
  assign T462 = ArrayRowModule_1_io_V_wire_en_5[4'he];
  assign T463 = ArrayRowModule_1_io_V_wire_en_5[4'hf];
  assign T464 = ArrayRowModule_1_io_V_wire_en_6[1'h0];
  assign T465 = ArrayRowModule_1_io_V_wire_en_6[1'h1];
  assign T466 = ArrayRowModule_1_io_V_wire_en_6[2'h2];
  assign T467 = ArrayRowModule_1_io_V_wire_en_6[2'h3];
  assign T468 = ArrayRowModule_1_io_V_wire_en_6[3'h4];
  assign T469 = ArrayRowModule_1_io_V_wire_en_6[3'h5];
  assign T470 = ArrayRowModule_1_io_V_wire_en_6[3'h6];
  assign T471 = ArrayRowModule_1_io_V_wire_en_6[3'h7];
  assign T472 = ArrayRowModule_1_io_V_wire_en_6[4'h8];
  assign T473 = ArrayRowModule_1_io_V_wire_en_6[4'h9];
  assign T474 = ArrayRowModule_1_io_V_wire_en_6[4'ha];
  assign T475 = ArrayRowModule_1_io_V_wire_en_6[4'hb];
  assign T476 = ArrayRowModule_1_io_V_wire_en_6[4'hc];
  assign T477 = ArrayRowModule_1_io_V_wire_en_6[4'hd];
  assign T478 = ArrayRowModule_1_io_V_wire_en_6[4'he];
  assign T479 = ArrayRowModule_1_io_V_wire_en_6[4'hf];
  assign T480 = ArrayRowModule_1_io_V_wire_en_7[1'h0];
  assign T481 = ArrayRowModule_1_io_V_wire_en_7[1'h1];
  assign T482 = ArrayRowModule_1_io_V_wire_en_7[2'h2];
  assign T483 = ArrayRowModule_1_io_V_wire_en_7[2'h3];
  assign T484 = ArrayRowModule_1_io_V_wire_en_7[3'h4];
  assign T485 = ArrayRowModule_1_io_V_wire_en_7[3'h5];
  assign T486 = ArrayRowModule_1_io_V_wire_en_7[3'h6];
  assign T487 = ArrayRowModule_1_io_V_wire_en_7[3'h7];
  assign T488 = ArrayRowModule_1_io_V_wire_en_7[4'h8];
  assign T489 = ArrayRowModule_1_io_V_wire_en_7[4'h9];
  assign T490 = ArrayRowModule_1_io_V_wire_en_7[4'ha];
  assign T491 = ArrayRowModule_1_io_V_wire_en_7[4'hb];
  assign T492 = ArrayRowModule_1_io_V_wire_en_7[4'hc];
  assign T493 = ArrayRowModule_1_io_V_wire_en_7[4'hd];
  assign T494 = ArrayRowModule_1_io_V_wire_en_7[4'he];
  assign T495 = ArrayRowModule_1_io_V_wire_en_7[4'hf];
  assign T496 = ArrayRowModule_1_io_V_wire_en_8[1'h0];
  assign T497 = ArrayRowModule_1_io_V_wire_en_8[1'h1];
  assign T498 = ArrayRowModule_1_io_V_wire_en_8[2'h2];
  assign T499 = ArrayRowModule_1_io_V_wire_en_8[2'h3];
  assign T500 = ArrayRowModule_1_io_V_wire_en_8[3'h4];
  assign T501 = ArrayRowModule_1_io_V_wire_en_8[3'h5];
  assign T502 = ArrayRowModule_1_io_V_wire_en_8[3'h6];
  assign T503 = ArrayRowModule_1_io_V_wire_en_8[3'h7];
  assign T504 = ArrayRowModule_1_io_V_wire_en_8[4'h8];
  assign T505 = ArrayRowModule_1_io_V_wire_en_8[4'h9];
  assign T506 = ArrayRowModule_1_io_V_wire_en_8[4'ha];
  assign T507 = ArrayRowModule_1_io_V_wire_en_8[4'hb];
  assign T508 = ArrayRowModule_1_io_V_wire_en_8[4'hc];
  assign T509 = ArrayRowModule_1_io_V_wire_en_8[4'hd];
  assign T510 = ArrayRowModule_1_io_V_wire_en_8[4'he];
  assign T511 = ArrayRowModule_1_io_V_wire_en_8[4'hf];
  assign T512 = ArrayRowModule_1_io_V_wire_en_9[1'h0];
  assign T513 = ArrayRowModule_1_io_V_wire_en_9[1'h1];
  assign T514 = ArrayRowModule_1_io_V_wire_en_9[2'h2];
  assign T515 = ArrayRowModule_1_io_V_wire_en_9[2'h3];
  assign T516 = ArrayRowModule_1_io_V_wire_en_9[3'h4];
  assign T517 = ArrayRowModule_1_io_V_wire_en_9[3'h5];
  assign T518 = ArrayRowModule_1_io_V_wire_en_9[3'h6];
  assign T519 = ArrayRowModule_1_io_V_wire_en_9[3'h7];
  assign T520 = ArrayRowModule_1_io_V_wire_en_9[4'h8];
  assign T521 = ArrayRowModule_1_io_V_wire_en_9[4'h9];
  assign T522 = ArrayRowModule_1_io_V_wire_en_9[4'ha];
  assign T523 = ArrayRowModule_1_io_V_wire_en_9[4'hb];
  assign T524 = ArrayRowModule_1_io_V_wire_en_9[4'hc];
  assign T525 = ArrayRowModule_1_io_V_wire_en_9[4'hd];
  assign T526 = ArrayRowModule_1_io_V_wire_en_9[4'he];
  assign T527 = ArrayRowModule_1_io_V_wire_en_9[4'hf];
  assign T528 = ArrayRowModule_1_io_V_wire_en_10[1'h0];
  assign T529 = ArrayRowModule_1_io_V_wire_en_10[1'h1];
  assign T530 = ArrayRowModule_1_io_V_wire_en_10[2'h2];
  assign T531 = ArrayRowModule_1_io_V_wire_en_10[2'h3];
  assign T532 = ArrayRowModule_1_io_V_wire_en_10[3'h4];
  assign T533 = ArrayRowModule_1_io_V_wire_en_10[3'h5];
  assign T534 = ArrayRowModule_1_io_V_wire_en_10[3'h6];
  assign T535 = ArrayRowModule_1_io_V_wire_en_10[3'h7];
  assign T536 = ArrayRowModule_1_io_V_wire_en_10[4'h8];
  assign T537 = ArrayRowModule_1_io_V_wire_en_10[4'h9];
  assign T538 = ArrayRowModule_1_io_V_wire_en_10[4'ha];
  assign T539 = ArrayRowModule_1_io_V_wire_en_10[4'hb];
  assign T540 = ArrayRowModule_1_io_V_wire_en_10[4'hc];
  assign T541 = ArrayRowModule_1_io_V_wire_en_10[4'hd];
  assign T542 = ArrayRowModule_1_io_V_wire_en_10[4'he];
  assign T543 = ArrayRowModule_1_io_V_wire_en_10[4'hf];
  assign T544 = ArrayRowModule_1_io_V_wire_en_11[1'h0];
  assign T545 = ArrayRowModule_1_io_V_wire_en_11[1'h1];
  assign T546 = ArrayRowModule_1_io_V_wire_en_11[2'h2];
  assign T547 = ArrayRowModule_1_io_V_wire_en_11[2'h3];
  assign T548 = ArrayRowModule_1_io_V_wire_en_11[3'h4];
  assign T549 = ArrayRowModule_1_io_V_wire_en_11[3'h5];
  assign T550 = ArrayRowModule_1_io_V_wire_en_11[3'h6];
  assign T551 = ArrayRowModule_1_io_V_wire_en_11[3'h7];
  assign T552 = ArrayRowModule_1_io_V_wire_en_11[4'h8];
  assign T553 = ArrayRowModule_1_io_V_wire_en_11[4'h9];
  assign T554 = ArrayRowModule_1_io_V_wire_en_11[4'ha];
  assign T555 = ArrayRowModule_1_io_V_wire_en_11[4'hb];
  assign T556 = ArrayRowModule_1_io_V_wire_en_11[4'hc];
  assign T557 = ArrayRowModule_1_io_V_wire_en_11[4'hd];
  assign T558 = ArrayRowModule_1_io_V_wire_en_11[4'he];
  assign T559 = ArrayRowModule_1_io_V_wire_en_11[4'hf];
  assign T560 = ArrayRowModule_1_io_V_wire_en_12[1'h0];
  assign T561 = ArrayRowModule_1_io_V_wire_en_12[1'h1];
  assign T562 = ArrayRowModule_1_io_V_wire_en_12[2'h2];
  assign T563 = ArrayRowModule_1_io_V_wire_en_12[2'h3];
  assign T564 = ArrayRowModule_1_io_V_wire_en_12[3'h4];
  assign T565 = ArrayRowModule_1_io_V_wire_en_12[3'h5];
  assign T566 = ArrayRowModule_1_io_V_wire_en_12[3'h6];
  assign T567 = ArrayRowModule_1_io_V_wire_en_12[3'h7];
  assign T568 = ArrayRowModule_1_io_V_wire_en_12[4'h8];
  assign T569 = ArrayRowModule_1_io_V_wire_en_12[4'h9];
  assign T570 = ArrayRowModule_1_io_V_wire_en_12[4'ha];
  assign T571 = ArrayRowModule_1_io_V_wire_en_12[4'hb];
  assign T572 = ArrayRowModule_1_io_V_wire_en_12[4'hc];
  assign T573 = ArrayRowModule_1_io_V_wire_en_12[4'hd];
  assign T574 = ArrayRowModule_1_io_V_wire_en_12[4'he];
  assign T575 = ArrayRowModule_1_io_V_wire_en_12[4'hf];
  assign T576 = ArrayRowModule_1_io_V_wire_en_13[1'h0];
  assign T577 = ArrayRowModule_1_io_V_wire_en_13[1'h1];
  assign T578 = ArrayRowModule_1_io_V_wire_en_13[2'h2];
  assign T579 = ArrayRowModule_1_io_V_wire_en_13[2'h3];
  assign T580 = ArrayRowModule_1_io_V_wire_en_13[3'h4];
  assign T581 = ArrayRowModule_1_io_V_wire_en_13[3'h5];
  assign T582 = ArrayRowModule_1_io_V_wire_en_13[3'h6];
  assign T583 = ArrayRowModule_1_io_V_wire_en_13[3'h7];
  assign T584 = ArrayRowModule_1_io_V_wire_en_13[4'h8];
  assign T585 = ArrayRowModule_1_io_V_wire_en_13[4'h9];
  assign T586 = ArrayRowModule_1_io_V_wire_en_13[4'ha];
  assign T587 = ArrayRowModule_1_io_V_wire_en_13[4'hb];
  assign T588 = ArrayRowModule_1_io_V_wire_en_13[4'hc];
  assign T589 = ArrayRowModule_1_io_V_wire_en_13[4'hd];
  assign T590 = ArrayRowModule_1_io_V_wire_en_13[4'he];
  assign T591 = ArrayRowModule_1_io_V_wire_en_13[4'hf];
  assign T592 = ArrayRowModule_1_io_V_wire_en_14[1'h0];
  assign T593 = ArrayRowModule_1_io_V_wire_en_14[1'h1];
  assign T594 = ArrayRowModule_1_io_V_wire_en_14[2'h2];
  assign T595 = ArrayRowModule_1_io_V_wire_en_14[2'h3];
  assign T596 = ArrayRowModule_1_io_V_wire_en_14[3'h4];
  assign T597 = ArrayRowModule_1_io_V_wire_en_14[3'h5];
  assign T598 = ArrayRowModule_1_io_V_wire_en_14[3'h6];
  assign T599 = ArrayRowModule_1_io_V_wire_en_14[3'h7];
  assign T600 = ArrayRowModule_1_io_V_wire_en_14[4'h8];
  assign T601 = ArrayRowModule_1_io_V_wire_en_14[4'h9];
  assign T602 = ArrayRowModule_1_io_V_wire_en_14[4'ha];
  assign T603 = ArrayRowModule_1_io_V_wire_en_14[4'hb];
  assign T604 = ArrayRowModule_1_io_V_wire_en_14[4'hc];
  assign T605 = ArrayRowModule_1_io_V_wire_en_14[4'hd];
  assign T606 = ArrayRowModule_1_io_V_wire_en_14[4'he];
  assign T607 = ArrayRowModule_1_io_V_wire_en_14[4'hf];
  assign T608 = ArrayRowModule_1_io_V_wire_en_15[1'h0];
  assign T609 = ArrayRowModule_1_io_V_wire_en_15[1'h1];
  assign T610 = ArrayRowModule_1_io_V_wire_en_15[2'h2];
  assign T611 = ArrayRowModule_1_io_V_wire_en_15[2'h3];
  assign T612 = ArrayRowModule_1_io_V_wire_en_15[3'h4];
  assign T613 = ArrayRowModule_1_io_V_wire_en_15[3'h5];
  assign T614 = ArrayRowModule_1_io_V_wire_en_15[3'h6];
  assign T615 = ArrayRowModule_1_io_V_wire_en_15[3'h7];
  assign T616 = ArrayRowModule_1_io_V_wire_en_15[4'h8];
  assign T617 = ArrayRowModule_1_io_V_wire_en_15[4'h9];
  assign T618 = ArrayRowModule_1_io_V_wire_en_15[4'ha];
  assign T619 = ArrayRowModule_1_io_V_wire_en_15[4'hb];
  assign T620 = ArrayRowModule_1_io_V_wire_en_15[4'hc];
  assign T621 = ArrayRowModule_1_io_V_wire_en_15[4'hd];
  assign T622 = ArrayRowModule_1_io_V_wire_en_15[4'he];
  assign T623 = ArrayRowModule_1_io_V_wire_en_15[4'hf];
  assign T624 = ArrayRowModule_1_io_V_wire_en_16[1'h0];
  assign T625 = ArrayRowModule_1_io_V_wire_en_16[1'h1];
  assign T626 = ArrayRowModule_1_io_V_wire_en_16[2'h2];
  assign T627 = ArrayRowModule_1_io_V_wire_en_16[2'h3];
  assign T628 = ArrayRowModule_1_io_V_wire_en_16[3'h4];
  assign T629 = ArrayRowModule_1_io_V_wire_en_16[3'h5];
  assign T630 = ArrayRowModule_1_io_V_wire_en_16[3'h6];
  assign T631 = ArrayRowModule_1_io_V_wire_en_16[3'h7];
  assign T632 = ArrayRowModule_1_io_V_wire_en_16[4'h8];
  assign T633 = ArrayRowModule_1_io_V_wire_en_16[4'h9];
  assign T634 = ArrayRowModule_1_io_V_wire_en_16[4'ha];
  assign T635 = ArrayRowModule_1_io_V_wire_en_16[4'hb];
  assign T636 = ArrayRowModule_1_io_V_wire_en_16[4'hc];
  assign T637 = ArrayRowModule_1_io_V_wire_en_16[4'hd];
  assign T638 = ArrayRowModule_1_io_V_wire_en_16[4'he];
  assign T639 = ArrayRowModule_1_io_V_wire_en_16[4'hf];
  assign T640 = ArrayRowModule_1_io_V_wire_en_17[1'h0];
  assign T641 = ArrayRowModule_1_io_V_wire_en_17[1'h1];
  assign T642 = ArrayRowModule_1_io_V_wire_en_17[2'h2];
  assign T643 = ArrayRowModule_1_io_V_wire_en_17[2'h3];
  assign T644 = ArrayRowModule_1_io_V_wire_en_17[3'h4];
  assign T645 = ArrayRowModule_1_io_V_wire_en_17[3'h5];
  assign T646 = ArrayRowModule_1_io_V_wire_en_17[3'h6];
  assign T647 = ArrayRowModule_1_io_V_wire_en_17[3'h7];
  assign T648 = ArrayRowModule_1_io_V_wire_en_17[4'h8];
  assign T649 = ArrayRowModule_1_io_V_wire_en_17[4'h9];
  assign T650 = ArrayRowModule_1_io_V_wire_en_17[4'ha];
  assign T651 = ArrayRowModule_1_io_V_wire_en_17[4'hb];
  assign T652 = ArrayRowModule_1_io_V_wire_en_17[4'hc];
  assign T653 = ArrayRowModule_1_io_V_wire_en_17[4'hd];
  assign T654 = ArrayRowModule_1_io_V_wire_en_17[4'he];
  assign T655 = ArrayRowModule_1_io_V_wire_en_17[4'hf];
  assign T656 = ArrayRowModule_1_io_V_wire_en_18[1'h0];
  assign T657 = ArrayRowModule_1_io_V_wire_en_18[1'h1];
  assign T658 = ArrayRowModule_1_io_V_wire_en_18[2'h2];
  assign T659 = ArrayRowModule_1_io_V_wire_en_18[2'h3];
  assign T660 = ArrayRowModule_1_io_V_wire_en_18[3'h4];
  assign T661 = ArrayRowModule_1_io_V_wire_en_18[3'h5];
  assign T662 = ArrayRowModule_1_io_V_wire_en_18[3'h6];
  assign T663 = ArrayRowModule_1_io_V_wire_en_18[3'h7];
  assign T664 = ArrayRowModule_1_io_V_wire_en_18[4'h8];
  assign T665 = ArrayRowModule_1_io_V_wire_en_18[4'h9];
  assign T666 = ArrayRowModule_1_io_V_wire_en_18[4'ha];
  assign T667 = ArrayRowModule_1_io_V_wire_en_18[4'hb];
  assign T668 = ArrayRowModule_1_io_V_wire_en_18[4'hc];
  assign T669 = ArrayRowModule_1_io_V_wire_en_18[4'hd];
  assign T670 = ArrayRowModule_1_io_V_wire_en_18[4'he];
  assign T671 = ArrayRowModule_1_io_V_wire_en_18[4'hf];
  assign T672 = ArrayRowModule_1_io_V_wire_en_19[1'h0];
  assign T673 = ArrayRowModule_1_io_V_wire_en_19[1'h1];
  assign T674 = ArrayRowModule_1_io_V_wire_en_19[2'h2];
  assign T675 = ArrayRowModule_1_io_V_wire_en_19[2'h3];
  assign T676 = ArrayRowModule_1_io_V_wire_en_19[3'h4];
  assign T677 = ArrayRowModule_1_io_V_wire_en_19[3'h5];
  assign T678 = ArrayRowModule_1_io_V_wire_en_19[3'h6];
  assign T679 = ArrayRowModule_1_io_V_wire_en_19[3'h7];
  assign T680 = ArrayRowModule_1_io_V_wire_en_19[4'h8];
  assign T681 = ArrayRowModule_1_io_V_wire_en_19[4'h9];
  assign T682 = ArrayRowModule_1_io_V_wire_en_19[4'ha];
  assign T683 = ArrayRowModule_1_io_V_wire_en_19[4'hb];
  assign T684 = ArrayRowModule_1_io_V_wire_en_19[4'hc];
  assign T685 = ArrayRowModule_1_io_V_wire_en_19[4'hd];
  assign T686 = ArrayRowModule_1_io_V_wire_en_19[4'he];
  assign T687 = ArrayRowModule_1_io_V_wire_en_19[4'hf];
  assign T688 = ArrayRowModule_1_io_V_wire_en_20[1'h0];
  assign T689 = ArrayRowModule_1_io_V_wire_en_20[1'h1];
  assign T690 = ArrayRowModule_1_io_V_wire_en_20[2'h2];
  assign T691 = ArrayRowModule_1_io_V_wire_en_20[2'h3];
  assign T692 = ArrayRowModule_1_io_V_wire_en_20[3'h4];
  assign T693 = ArrayRowModule_1_io_V_wire_en_20[3'h5];
  assign T694 = ArrayRowModule_1_io_V_wire_en_20[3'h6];
  assign T695 = ArrayRowModule_1_io_V_wire_en_20[3'h7];
  assign T696 = ArrayRowModule_1_io_V_wire_en_20[4'h8];
  assign T697 = ArrayRowModule_1_io_V_wire_en_20[4'h9];
  assign T698 = ArrayRowModule_1_io_V_wire_en_20[4'ha];
  assign T699 = ArrayRowModule_1_io_V_wire_en_20[4'hb];
  assign T700 = ArrayRowModule_1_io_V_wire_en_20[4'hc];
  assign T701 = ArrayRowModule_1_io_V_wire_en_20[4'hd];
  assign T702 = ArrayRowModule_1_io_V_wire_en_20[4'he];
  assign T703 = ArrayRowModule_1_io_V_wire_en_20[4'hf];
  assign T704 = ArrayRowModule_1_io_V_wire_en_21[1'h0];
  assign T705 = ArrayRowModule_1_io_V_wire_en_21[1'h1];
  assign T706 = ArrayRowModule_1_io_V_wire_en_21[2'h2];
  assign T707 = ArrayRowModule_1_io_V_wire_en_21[2'h3];
  assign T708 = ArrayRowModule_1_io_V_wire_en_21[3'h4];
  assign T709 = ArrayRowModule_1_io_V_wire_en_21[3'h5];
  assign T710 = ArrayRowModule_1_io_V_wire_en_21[3'h6];
  assign T711 = ArrayRowModule_1_io_V_wire_en_21[3'h7];
  assign T712 = ArrayRowModule_1_io_V_wire_en_21[4'h8];
  assign T713 = ArrayRowModule_1_io_V_wire_en_21[4'h9];
  assign T714 = ArrayRowModule_1_io_V_wire_en_21[4'ha];
  assign T715 = ArrayRowModule_1_io_V_wire_en_21[4'hb];
  assign T716 = ArrayRowModule_1_io_V_wire_en_21[4'hc];
  assign T717 = ArrayRowModule_1_io_V_wire_en_21[4'hd];
  assign T718 = ArrayRowModule_1_io_V_wire_en_21[4'he];
  assign T719 = ArrayRowModule_1_io_V_wire_en_21[4'hf];
  assign T720 = ArrayRowModule_1_io_V_wire_en_22[1'h0];
  assign T721 = ArrayRowModule_1_io_V_wire_en_22[1'h1];
  assign T722 = ArrayRowModule_1_io_V_wire_en_22[2'h2];
  assign T723 = ArrayRowModule_1_io_V_wire_en_22[2'h3];
  assign T724 = ArrayRowModule_1_io_V_wire_en_22[3'h4];
  assign T725 = ArrayRowModule_1_io_V_wire_en_22[3'h5];
  assign T726 = ArrayRowModule_1_io_V_wire_en_22[3'h6];
  assign T727 = ArrayRowModule_1_io_V_wire_en_22[3'h7];
  assign T728 = ArrayRowModule_1_io_V_wire_en_22[4'h8];
  assign T729 = ArrayRowModule_1_io_V_wire_en_22[4'h9];
  assign T730 = ArrayRowModule_1_io_V_wire_en_22[4'ha];
  assign T731 = ArrayRowModule_1_io_V_wire_en_22[4'hb];
  assign T732 = ArrayRowModule_1_io_V_wire_en_22[4'hc];
  assign T733 = ArrayRowModule_1_io_V_wire_en_22[4'hd];
  assign T734 = ArrayRowModule_1_io_V_wire_en_22[4'he];
  assign T735 = ArrayRowModule_1_io_V_wire_en_22[4'hf];
  assign T736 = ArrayRowModule_2_io_V_wire_en_0[1'h0];
  assign T737 = ArrayRowModule_2_io_V_wire_en_0[1'h1];
  assign T738 = ArrayRowModule_2_io_V_wire_en_0[2'h2];
  assign T739 = ArrayRowModule_2_io_V_wire_en_0[2'h3];
  assign T740 = ArrayRowModule_2_io_V_wire_en_0[3'h4];
  assign T741 = ArrayRowModule_2_io_V_wire_en_0[3'h5];
  assign T742 = ArrayRowModule_2_io_V_wire_en_0[3'h6];
  assign T743 = ArrayRowModule_2_io_V_wire_en_0[3'h7];
  assign T744 = ArrayRowModule_2_io_V_wire_en_0[4'h8];
  assign T745 = ArrayRowModule_2_io_V_wire_en_0[4'h9];
  assign T746 = ArrayRowModule_2_io_V_wire_en_0[4'ha];
  assign T747 = ArrayRowModule_2_io_V_wire_en_0[4'hb];
  assign T748 = ArrayRowModule_2_io_V_wire_en_0[4'hc];
  assign T749 = ArrayRowModule_2_io_V_wire_en_0[4'hd];
  assign T750 = ArrayRowModule_2_io_V_wire_en_0[4'he];
  assign T751 = ArrayRowModule_2_io_V_wire_en_0[4'hf];
  assign T752 = ArrayRowModule_2_io_V_wire_en_1[1'h0];
  assign T753 = ArrayRowModule_2_io_V_wire_en_1[1'h1];
  assign T754 = ArrayRowModule_2_io_V_wire_en_1[2'h2];
  assign T755 = ArrayRowModule_2_io_V_wire_en_1[2'h3];
  assign T756 = ArrayRowModule_2_io_V_wire_en_1[3'h4];
  assign T757 = ArrayRowModule_2_io_V_wire_en_1[3'h5];
  assign T758 = ArrayRowModule_2_io_V_wire_en_1[3'h6];
  assign T759 = ArrayRowModule_2_io_V_wire_en_1[3'h7];
  assign T760 = ArrayRowModule_2_io_V_wire_en_1[4'h8];
  assign T761 = ArrayRowModule_2_io_V_wire_en_1[4'h9];
  assign T762 = ArrayRowModule_2_io_V_wire_en_1[4'ha];
  assign T763 = ArrayRowModule_2_io_V_wire_en_1[4'hb];
  assign T764 = ArrayRowModule_2_io_V_wire_en_1[4'hc];
  assign T765 = ArrayRowModule_2_io_V_wire_en_1[4'hd];
  assign T766 = ArrayRowModule_2_io_V_wire_en_1[4'he];
  assign T767 = ArrayRowModule_2_io_V_wire_en_1[4'hf];
  assign T768 = ArrayRowModule_2_io_V_wire_en_2[1'h0];
  assign T769 = ArrayRowModule_2_io_V_wire_en_2[1'h1];
  assign T770 = ArrayRowModule_2_io_V_wire_en_2[2'h2];
  assign T771 = ArrayRowModule_2_io_V_wire_en_2[2'h3];
  assign T772 = ArrayRowModule_2_io_V_wire_en_2[3'h4];
  assign T773 = ArrayRowModule_2_io_V_wire_en_2[3'h5];
  assign T774 = ArrayRowModule_2_io_V_wire_en_2[3'h6];
  assign T775 = ArrayRowModule_2_io_V_wire_en_2[3'h7];
  assign T776 = ArrayRowModule_2_io_V_wire_en_2[4'h8];
  assign T777 = ArrayRowModule_2_io_V_wire_en_2[4'h9];
  assign T778 = ArrayRowModule_2_io_V_wire_en_2[4'ha];
  assign T779 = ArrayRowModule_2_io_V_wire_en_2[4'hb];
  assign T780 = ArrayRowModule_2_io_V_wire_en_2[4'hc];
  assign T781 = ArrayRowModule_2_io_V_wire_en_2[4'hd];
  assign T782 = ArrayRowModule_2_io_V_wire_en_2[4'he];
  assign T783 = ArrayRowModule_2_io_V_wire_en_2[4'hf];
  assign T784 = ArrayRowModule_2_io_V_wire_en_3[1'h0];
  assign T785 = ArrayRowModule_2_io_V_wire_en_3[1'h1];
  assign T786 = ArrayRowModule_2_io_V_wire_en_3[2'h2];
  assign T787 = ArrayRowModule_2_io_V_wire_en_3[2'h3];
  assign T788 = ArrayRowModule_2_io_V_wire_en_3[3'h4];
  assign T789 = ArrayRowModule_2_io_V_wire_en_3[3'h5];
  assign T790 = ArrayRowModule_2_io_V_wire_en_3[3'h6];
  assign T791 = ArrayRowModule_2_io_V_wire_en_3[3'h7];
  assign T792 = ArrayRowModule_2_io_V_wire_en_3[4'h8];
  assign T793 = ArrayRowModule_2_io_V_wire_en_3[4'h9];
  assign T794 = ArrayRowModule_2_io_V_wire_en_3[4'ha];
  assign T795 = ArrayRowModule_2_io_V_wire_en_3[4'hb];
  assign T796 = ArrayRowModule_2_io_V_wire_en_3[4'hc];
  assign T797 = ArrayRowModule_2_io_V_wire_en_3[4'hd];
  assign T798 = ArrayRowModule_2_io_V_wire_en_3[4'he];
  assign T799 = ArrayRowModule_2_io_V_wire_en_3[4'hf];
  assign T800 = ArrayRowModule_2_io_V_wire_en_4[1'h0];
  assign T801 = ArrayRowModule_2_io_V_wire_en_4[1'h1];
  assign T802 = ArrayRowModule_2_io_V_wire_en_4[2'h2];
  assign T803 = ArrayRowModule_2_io_V_wire_en_4[2'h3];
  assign T804 = ArrayRowModule_2_io_V_wire_en_4[3'h4];
  assign T805 = ArrayRowModule_2_io_V_wire_en_4[3'h5];
  assign T806 = ArrayRowModule_2_io_V_wire_en_4[3'h6];
  assign T807 = ArrayRowModule_2_io_V_wire_en_4[3'h7];
  assign T808 = ArrayRowModule_2_io_V_wire_en_4[4'h8];
  assign T809 = ArrayRowModule_2_io_V_wire_en_4[4'h9];
  assign T810 = ArrayRowModule_2_io_V_wire_en_4[4'ha];
  assign T811 = ArrayRowModule_2_io_V_wire_en_4[4'hb];
  assign T812 = ArrayRowModule_2_io_V_wire_en_4[4'hc];
  assign T813 = ArrayRowModule_2_io_V_wire_en_4[4'hd];
  assign T814 = ArrayRowModule_2_io_V_wire_en_4[4'he];
  assign T815 = ArrayRowModule_2_io_V_wire_en_4[4'hf];
  assign T816 = ArrayRowModule_2_io_V_wire_en_5[1'h0];
  assign T817 = ArrayRowModule_2_io_V_wire_en_5[1'h1];
  assign T818 = ArrayRowModule_2_io_V_wire_en_5[2'h2];
  assign T819 = ArrayRowModule_2_io_V_wire_en_5[2'h3];
  assign T820 = ArrayRowModule_2_io_V_wire_en_5[3'h4];
  assign T821 = ArrayRowModule_2_io_V_wire_en_5[3'h5];
  assign T822 = ArrayRowModule_2_io_V_wire_en_5[3'h6];
  assign T823 = ArrayRowModule_2_io_V_wire_en_5[3'h7];
  assign T824 = ArrayRowModule_2_io_V_wire_en_5[4'h8];
  assign T825 = ArrayRowModule_2_io_V_wire_en_5[4'h9];
  assign T826 = ArrayRowModule_2_io_V_wire_en_5[4'ha];
  assign T827 = ArrayRowModule_2_io_V_wire_en_5[4'hb];
  assign T828 = ArrayRowModule_2_io_V_wire_en_5[4'hc];
  assign T829 = ArrayRowModule_2_io_V_wire_en_5[4'hd];
  assign T830 = ArrayRowModule_2_io_V_wire_en_5[4'he];
  assign T831 = ArrayRowModule_2_io_V_wire_en_5[4'hf];
  assign T832 = ArrayRowModule_2_io_V_wire_en_6[1'h0];
  assign T833 = ArrayRowModule_2_io_V_wire_en_6[1'h1];
  assign T834 = ArrayRowModule_2_io_V_wire_en_6[2'h2];
  assign T835 = ArrayRowModule_2_io_V_wire_en_6[2'h3];
  assign T836 = ArrayRowModule_2_io_V_wire_en_6[3'h4];
  assign T837 = ArrayRowModule_2_io_V_wire_en_6[3'h5];
  assign T838 = ArrayRowModule_2_io_V_wire_en_6[3'h6];
  assign T839 = ArrayRowModule_2_io_V_wire_en_6[3'h7];
  assign T840 = ArrayRowModule_2_io_V_wire_en_6[4'h8];
  assign T841 = ArrayRowModule_2_io_V_wire_en_6[4'h9];
  assign T842 = ArrayRowModule_2_io_V_wire_en_6[4'ha];
  assign T843 = ArrayRowModule_2_io_V_wire_en_6[4'hb];
  assign T844 = ArrayRowModule_2_io_V_wire_en_6[4'hc];
  assign T845 = ArrayRowModule_2_io_V_wire_en_6[4'hd];
  assign T846 = ArrayRowModule_2_io_V_wire_en_6[4'he];
  assign T847 = ArrayRowModule_2_io_V_wire_en_6[4'hf];
  assign T848 = ArrayRowModule_2_io_V_wire_en_7[1'h0];
  assign T849 = ArrayRowModule_2_io_V_wire_en_7[1'h1];
  assign T850 = ArrayRowModule_2_io_V_wire_en_7[2'h2];
  assign T851 = ArrayRowModule_2_io_V_wire_en_7[2'h3];
  assign T852 = ArrayRowModule_2_io_V_wire_en_7[3'h4];
  assign T853 = ArrayRowModule_2_io_V_wire_en_7[3'h5];
  assign T854 = ArrayRowModule_2_io_V_wire_en_7[3'h6];
  assign T855 = ArrayRowModule_2_io_V_wire_en_7[3'h7];
  assign T856 = ArrayRowModule_2_io_V_wire_en_7[4'h8];
  assign T857 = ArrayRowModule_2_io_V_wire_en_7[4'h9];
  assign T858 = ArrayRowModule_2_io_V_wire_en_7[4'ha];
  assign T859 = ArrayRowModule_2_io_V_wire_en_7[4'hb];
  assign T860 = ArrayRowModule_2_io_V_wire_en_7[4'hc];
  assign T861 = ArrayRowModule_2_io_V_wire_en_7[4'hd];
  assign T862 = ArrayRowModule_2_io_V_wire_en_7[4'he];
  assign T863 = ArrayRowModule_2_io_V_wire_en_7[4'hf];
  assign T864 = ArrayRowModule_2_io_V_wire_en_8[1'h0];
  assign T865 = ArrayRowModule_2_io_V_wire_en_8[1'h1];
  assign T866 = ArrayRowModule_2_io_V_wire_en_8[2'h2];
  assign T867 = ArrayRowModule_2_io_V_wire_en_8[2'h3];
  assign T868 = ArrayRowModule_2_io_V_wire_en_8[3'h4];
  assign T869 = ArrayRowModule_2_io_V_wire_en_8[3'h5];
  assign T870 = ArrayRowModule_2_io_V_wire_en_8[3'h6];
  assign T871 = ArrayRowModule_2_io_V_wire_en_8[3'h7];
  assign T872 = ArrayRowModule_2_io_V_wire_en_8[4'h8];
  assign T873 = ArrayRowModule_2_io_V_wire_en_8[4'h9];
  assign T874 = ArrayRowModule_2_io_V_wire_en_8[4'ha];
  assign T875 = ArrayRowModule_2_io_V_wire_en_8[4'hb];
  assign T876 = ArrayRowModule_2_io_V_wire_en_8[4'hc];
  assign T877 = ArrayRowModule_2_io_V_wire_en_8[4'hd];
  assign T878 = ArrayRowModule_2_io_V_wire_en_8[4'he];
  assign T879 = ArrayRowModule_2_io_V_wire_en_8[4'hf];
  assign T880 = ArrayRowModule_2_io_V_wire_en_9[1'h0];
  assign T881 = ArrayRowModule_2_io_V_wire_en_9[1'h1];
  assign T882 = ArrayRowModule_2_io_V_wire_en_9[2'h2];
  assign T883 = ArrayRowModule_2_io_V_wire_en_9[2'h3];
  assign T884 = ArrayRowModule_2_io_V_wire_en_9[3'h4];
  assign T885 = ArrayRowModule_2_io_V_wire_en_9[3'h5];
  assign T886 = ArrayRowModule_2_io_V_wire_en_9[3'h6];
  assign T887 = ArrayRowModule_2_io_V_wire_en_9[3'h7];
  assign T888 = ArrayRowModule_2_io_V_wire_en_9[4'h8];
  assign T889 = ArrayRowModule_2_io_V_wire_en_9[4'h9];
  assign T890 = ArrayRowModule_2_io_V_wire_en_9[4'ha];
  assign T891 = ArrayRowModule_2_io_V_wire_en_9[4'hb];
  assign T892 = ArrayRowModule_2_io_V_wire_en_9[4'hc];
  assign T893 = ArrayRowModule_2_io_V_wire_en_9[4'hd];
  assign T894 = ArrayRowModule_2_io_V_wire_en_9[4'he];
  assign T895 = ArrayRowModule_2_io_V_wire_en_9[4'hf];
  assign T896 = ArrayRowModule_2_io_V_wire_en_10[1'h0];
  assign T897 = ArrayRowModule_2_io_V_wire_en_10[1'h1];
  assign T898 = ArrayRowModule_2_io_V_wire_en_10[2'h2];
  assign T899 = ArrayRowModule_2_io_V_wire_en_10[2'h3];
  assign T900 = ArrayRowModule_2_io_V_wire_en_10[3'h4];
  assign T901 = ArrayRowModule_2_io_V_wire_en_10[3'h5];
  assign T902 = ArrayRowModule_2_io_V_wire_en_10[3'h6];
  assign T903 = ArrayRowModule_2_io_V_wire_en_10[3'h7];
  assign T904 = ArrayRowModule_2_io_V_wire_en_10[4'h8];
  assign T905 = ArrayRowModule_2_io_V_wire_en_10[4'h9];
  assign T906 = ArrayRowModule_2_io_V_wire_en_10[4'ha];
  assign T907 = ArrayRowModule_2_io_V_wire_en_10[4'hb];
  assign T908 = ArrayRowModule_2_io_V_wire_en_10[4'hc];
  assign T909 = ArrayRowModule_2_io_V_wire_en_10[4'hd];
  assign T910 = ArrayRowModule_2_io_V_wire_en_10[4'he];
  assign T911 = ArrayRowModule_2_io_V_wire_en_10[4'hf];
  assign T912 = ArrayRowModule_2_io_V_wire_en_11[1'h0];
  assign T913 = ArrayRowModule_2_io_V_wire_en_11[1'h1];
  assign T914 = ArrayRowModule_2_io_V_wire_en_11[2'h2];
  assign T915 = ArrayRowModule_2_io_V_wire_en_11[2'h3];
  assign T916 = ArrayRowModule_2_io_V_wire_en_11[3'h4];
  assign T917 = ArrayRowModule_2_io_V_wire_en_11[3'h5];
  assign T918 = ArrayRowModule_2_io_V_wire_en_11[3'h6];
  assign T919 = ArrayRowModule_2_io_V_wire_en_11[3'h7];
  assign T920 = ArrayRowModule_2_io_V_wire_en_11[4'h8];
  assign T921 = ArrayRowModule_2_io_V_wire_en_11[4'h9];
  assign T922 = ArrayRowModule_2_io_V_wire_en_11[4'ha];
  assign T923 = ArrayRowModule_2_io_V_wire_en_11[4'hb];
  assign T924 = ArrayRowModule_2_io_V_wire_en_11[4'hc];
  assign T925 = ArrayRowModule_2_io_V_wire_en_11[4'hd];
  assign T926 = ArrayRowModule_2_io_V_wire_en_11[4'he];
  assign T927 = ArrayRowModule_2_io_V_wire_en_11[4'hf];
  assign T928 = ArrayRowModule_2_io_V_wire_en_12[1'h0];
  assign T929 = ArrayRowModule_2_io_V_wire_en_12[1'h1];
  assign T930 = ArrayRowModule_2_io_V_wire_en_12[2'h2];
  assign T931 = ArrayRowModule_2_io_V_wire_en_12[2'h3];
  assign T932 = ArrayRowModule_2_io_V_wire_en_12[3'h4];
  assign T933 = ArrayRowModule_2_io_V_wire_en_12[3'h5];
  assign T934 = ArrayRowModule_2_io_V_wire_en_12[3'h6];
  assign T935 = ArrayRowModule_2_io_V_wire_en_12[3'h7];
  assign T936 = ArrayRowModule_2_io_V_wire_en_12[4'h8];
  assign T937 = ArrayRowModule_2_io_V_wire_en_12[4'h9];
  assign T938 = ArrayRowModule_2_io_V_wire_en_12[4'ha];
  assign T939 = ArrayRowModule_2_io_V_wire_en_12[4'hb];
  assign T940 = ArrayRowModule_2_io_V_wire_en_12[4'hc];
  assign T941 = ArrayRowModule_2_io_V_wire_en_12[4'hd];
  assign T942 = ArrayRowModule_2_io_V_wire_en_12[4'he];
  assign T943 = ArrayRowModule_2_io_V_wire_en_12[4'hf];
  assign T944 = ArrayRowModule_2_io_V_wire_en_13[1'h0];
  assign T945 = ArrayRowModule_2_io_V_wire_en_13[1'h1];
  assign T946 = ArrayRowModule_2_io_V_wire_en_13[2'h2];
  assign T947 = ArrayRowModule_2_io_V_wire_en_13[2'h3];
  assign T948 = ArrayRowModule_2_io_V_wire_en_13[3'h4];
  assign T949 = ArrayRowModule_2_io_V_wire_en_13[3'h5];
  assign T950 = ArrayRowModule_2_io_V_wire_en_13[3'h6];
  assign T951 = ArrayRowModule_2_io_V_wire_en_13[3'h7];
  assign T952 = ArrayRowModule_2_io_V_wire_en_13[4'h8];
  assign T953 = ArrayRowModule_2_io_V_wire_en_13[4'h9];
  assign T954 = ArrayRowModule_2_io_V_wire_en_13[4'ha];
  assign T955 = ArrayRowModule_2_io_V_wire_en_13[4'hb];
  assign T956 = ArrayRowModule_2_io_V_wire_en_13[4'hc];
  assign T957 = ArrayRowModule_2_io_V_wire_en_13[4'hd];
  assign T958 = ArrayRowModule_2_io_V_wire_en_13[4'he];
  assign T959 = ArrayRowModule_2_io_V_wire_en_13[4'hf];
  assign T960 = ArrayRowModule_2_io_V_wire_en_14[1'h0];
  assign T961 = ArrayRowModule_2_io_V_wire_en_14[1'h1];
  assign T962 = ArrayRowModule_2_io_V_wire_en_14[2'h2];
  assign T963 = ArrayRowModule_2_io_V_wire_en_14[2'h3];
  assign T964 = ArrayRowModule_2_io_V_wire_en_14[3'h4];
  assign T965 = ArrayRowModule_2_io_V_wire_en_14[3'h5];
  assign T966 = ArrayRowModule_2_io_V_wire_en_14[3'h6];
  assign T967 = ArrayRowModule_2_io_V_wire_en_14[3'h7];
  assign T968 = ArrayRowModule_2_io_V_wire_en_14[4'h8];
  assign T969 = ArrayRowModule_2_io_V_wire_en_14[4'h9];
  assign T970 = ArrayRowModule_2_io_V_wire_en_14[4'ha];
  assign T971 = ArrayRowModule_2_io_V_wire_en_14[4'hb];
  assign T972 = ArrayRowModule_2_io_V_wire_en_14[4'hc];
  assign T973 = ArrayRowModule_2_io_V_wire_en_14[4'hd];
  assign T974 = ArrayRowModule_2_io_V_wire_en_14[4'he];
  assign T975 = ArrayRowModule_2_io_V_wire_en_14[4'hf];
  assign T976 = ArrayRowModule_2_io_V_wire_en_15[1'h0];
  assign T977 = ArrayRowModule_2_io_V_wire_en_15[1'h1];
  assign T978 = ArrayRowModule_2_io_V_wire_en_15[2'h2];
  assign T979 = ArrayRowModule_2_io_V_wire_en_15[2'h3];
  assign T980 = ArrayRowModule_2_io_V_wire_en_15[3'h4];
  assign T981 = ArrayRowModule_2_io_V_wire_en_15[3'h5];
  assign T982 = ArrayRowModule_2_io_V_wire_en_15[3'h6];
  assign T983 = ArrayRowModule_2_io_V_wire_en_15[3'h7];
  assign T984 = ArrayRowModule_2_io_V_wire_en_15[4'h8];
  assign T985 = ArrayRowModule_2_io_V_wire_en_15[4'h9];
  assign T986 = ArrayRowModule_2_io_V_wire_en_15[4'ha];
  assign T987 = ArrayRowModule_2_io_V_wire_en_15[4'hb];
  assign T988 = ArrayRowModule_2_io_V_wire_en_15[4'hc];
  assign T989 = ArrayRowModule_2_io_V_wire_en_15[4'hd];
  assign T990 = ArrayRowModule_2_io_V_wire_en_15[4'he];
  assign T991 = ArrayRowModule_2_io_V_wire_en_15[4'hf];
  assign T992 = ArrayRowModule_2_io_V_wire_en_16[1'h0];
  assign T993 = ArrayRowModule_2_io_V_wire_en_16[1'h1];
  assign T994 = ArrayRowModule_2_io_V_wire_en_16[2'h2];
  assign T995 = ArrayRowModule_2_io_V_wire_en_16[2'h3];
  assign T996 = ArrayRowModule_2_io_V_wire_en_16[3'h4];
  assign T997 = ArrayRowModule_2_io_V_wire_en_16[3'h5];
  assign T998 = ArrayRowModule_2_io_V_wire_en_16[3'h6];
  assign T999 = ArrayRowModule_2_io_V_wire_en_16[3'h7];
  assign T1000 = ArrayRowModule_2_io_V_wire_en_16[4'h8];
  assign T1001 = ArrayRowModule_2_io_V_wire_en_16[4'h9];
  assign T1002 = ArrayRowModule_2_io_V_wire_en_16[4'ha];
  assign T1003 = ArrayRowModule_2_io_V_wire_en_16[4'hb];
  assign T1004 = ArrayRowModule_2_io_V_wire_en_16[4'hc];
  assign T1005 = ArrayRowModule_2_io_V_wire_en_16[4'hd];
  assign T1006 = ArrayRowModule_2_io_V_wire_en_16[4'he];
  assign T1007 = ArrayRowModule_2_io_V_wire_en_16[4'hf];
  assign T1008 = ArrayRowModule_2_io_V_wire_en_17[1'h0];
  assign T1009 = ArrayRowModule_2_io_V_wire_en_17[1'h1];
  assign T1010 = ArrayRowModule_2_io_V_wire_en_17[2'h2];
  assign T1011 = ArrayRowModule_2_io_V_wire_en_17[2'h3];
  assign T1012 = ArrayRowModule_2_io_V_wire_en_17[3'h4];
  assign T1013 = ArrayRowModule_2_io_V_wire_en_17[3'h5];
  assign T1014 = ArrayRowModule_2_io_V_wire_en_17[3'h6];
  assign T1015 = ArrayRowModule_2_io_V_wire_en_17[3'h7];
  assign T1016 = ArrayRowModule_2_io_V_wire_en_17[4'h8];
  assign T1017 = ArrayRowModule_2_io_V_wire_en_17[4'h9];
  assign T1018 = ArrayRowModule_2_io_V_wire_en_17[4'ha];
  assign T1019 = ArrayRowModule_2_io_V_wire_en_17[4'hb];
  assign T1020 = ArrayRowModule_2_io_V_wire_en_17[4'hc];
  assign T1021 = ArrayRowModule_2_io_V_wire_en_17[4'hd];
  assign T1022 = ArrayRowModule_2_io_V_wire_en_17[4'he];
  assign T1023 = ArrayRowModule_2_io_V_wire_en_17[4'hf];
  assign T1024 = ArrayRowModule_2_io_V_wire_en_18[1'h0];
  assign T1025 = ArrayRowModule_2_io_V_wire_en_18[1'h1];
  assign T1026 = ArrayRowModule_2_io_V_wire_en_18[2'h2];
  assign T1027 = ArrayRowModule_2_io_V_wire_en_18[2'h3];
  assign T1028 = ArrayRowModule_2_io_V_wire_en_18[3'h4];
  assign T1029 = ArrayRowModule_2_io_V_wire_en_18[3'h5];
  assign T1030 = ArrayRowModule_2_io_V_wire_en_18[3'h6];
  assign T1031 = ArrayRowModule_2_io_V_wire_en_18[3'h7];
  assign T1032 = ArrayRowModule_2_io_V_wire_en_18[4'h8];
  assign T1033 = ArrayRowModule_2_io_V_wire_en_18[4'h9];
  assign T1034 = ArrayRowModule_2_io_V_wire_en_18[4'ha];
  assign T1035 = ArrayRowModule_2_io_V_wire_en_18[4'hb];
  assign T1036 = ArrayRowModule_2_io_V_wire_en_18[4'hc];
  assign T1037 = ArrayRowModule_2_io_V_wire_en_18[4'hd];
  assign T1038 = ArrayRowModule_2_io_V_wire_en_18[4'he];
  assign T1039 = ArrayRowModule_2_io_V_wire_en_18[4'hf];
  assign T1040 = ArrayRowModule_2_io_V_wire_en_19[1'h0];
  assign T1041 = ArrayRowModule_2_io_V_wire_en_19[1'h1];
  assign T1042 = ArrayRowModule_2_io_V_wire_en_19[2'h2];
  assign T1043 = ArrayRowModule_2_io_V_wire_en_19[2'h3];
  assign T1044 = ArrayRowModule_2_io_V_wire_en_19[3'h4];
  assign T1045 = ArrayRowModule_2_io_V_wire_en_19[3'h5];
  assign T1046 = ArrayRowModule_2_io_V_wire_en_19[3'h6];
  assign T1047 = ArrayRowModule_2_io_V_wire_en_19[3'h7];
  assign T1048 = ArrayRowModule_2_io_V_wire_en_19[4'h8];
  assign T1049 = ArrayRowModule_2_io_V_wire_en_19[4'h9];
  assign T1050 = ArrayRowModule_2_io_V_wire_en_19[4'ha];
  assign T1051 = ArrayRowModule_2_io_V_wire_en_19[4'hb];
  assign T1052 = ArrayRowModule_2_io_V_wire_en_19[4'hc];
  assign T1053 = ArrayRowModule_2_io_V_wire_en_19[4'hd];
  assign T1054 = ArrayRowModule_2_io_V_wire_en_19[4'he];
  assign T1055 = ArrayRowModule_2_io_V_wire_en_19[4'hf];
  assign T1056 = ArrayRowModule_2_io_V_wire_en_20[1'h0];
  assign T1057 = ArrayRowModule_2_io_V_wire_en_20[1'h1];
  assign T1058 = ArrayRowModule_2_io_V_wire_en_20[2'h2];
  assign T1059 = ArrayRowModule_2_io_V_wire_en_20[2'h3];
  assign T1060 = ArrayRowModule_2_io_V_wire_en_20[3'h4];
  assign T1061 = ArrayRowModule_2_io_V_wire_en_20[3'h5];
  assign T1062 = ArrayRowModule_2_io_V_wire_en_20[3'h6];
  assign T1063 = ArrayRowModule_2_io_V_wire_en_20[3'h7];
  assign T1064 = ArrayRowModule_2_io_V_wire_en_20[4'h8];
  assign T1065 = ArrayRowModule_2_io_V_wire_en_20[4'h9];
  assign T1066 = ArrayRowModule_2_io_V_wire_en_20[4'ha];
  assign T1067 = ArrayRowModule_2_io_V_wire_en_20[4'hb];
  assign T1068 = ArrayRowModule_2_io_V_wire_en_20[4'hc];
  assign T1069 = ArrayRowModule_2_io_V_wire_en_20[4'hd];
  assign T1070 = ArrayRowModule_2_io_V_wire_en_20[4'he];
  assign T1071 = ArrayRowModule_2_io_V_wire_en_20[4'hf];
  assign T1072 = ArrayRowModule_2_io_V_wire_en_21[1'h0];
  assign T1073 = ArrayRowModule_2_io_V_wire_en_21[1'h1];
  assign T1074 = ArrayRowModule_2_io_V_wire_en_21[2'h2];
  assign T1075 = ArrayRowModule_2_io_V_wire_en_21[2'h3];
  assign T1076 = ArrayRowModule_2_io_V_wire_en_21[3'h4];
  assign T1077 = ArrayRowModule_2_io_V_wire_en_21[3'h5];
  assign T1078 = ArrayRowModule_2_io_V_wire_en_21[3'h6];
  assign T1079 = ArrayRowModule_2_io_V_wire_en_21[3'h7];
  assign T1080 = ArrayRowModule_2_io_V_wire_en_21[4'h8];
  assign T1081 = ArrayRowModule_2_io_V_wire_en_21[4'h9];
  assign T1082 = ArrayRowModule_2_io_V_wire_en_21[4'ha];
  assign T1083 = ArrayRowModule_2_io_V_wire_en_21[4'hb];
  assign T1084 = ArrayRowModule_2_io_V_wire_en_21[4'hc];
  assign T1085 = ArrayRowModule_2_io_V_wire_en_21[4'hd];
  assign T1086 = ArrayRowModule_2_io_V_wire_en_21[4'he];
  assign T1087 = ArrayRowModule_2_io_V_wire_en_21[4'hf];
  assign T1088 = ArrayRowModule_2_io_V_wire_en_22[1'h0];
  assign T1089 = ArrayRowModule_2_io_V_wire_en_22[1'h1];
  assign T1090 = ArrayRowModule_2_io_V_wire_en_22[2'h2];
  assign T1091 = ArrayRowModule_2_io_V_wire_en_22[2'h3];
  assign T1092 = ArrayRowModule_2_io_V_wire_en_22[3'h4];
  assign T1093 = ArrayRowModule_2_io_V_wire_en_22[3'h5];
  assign T1094 = ArrayRowModule_2_io_V_wire_en_22[3'h6];
  assign T1095 = ArrayRowModule_2_io_V_wire_en_22[3'h7];
  assign T1096 = ArrayRowModule_2_io_V_wire_en_22[4'h8];
  assign T1097 = ArrayRowModule_2_io_V_wire_en_22[4'h9];
  assign T1098 = ArrayRowModule_2_io_V_wire_en_22[4'ha];
  assign T1099 = ArrayRowModule_2_io_V_wire_en_22[4'hb];
  assign T1100 = ArrayRowModule_2_io_V_wire_en_22[4'hc];
  assign T1101 = ArrayRowModule_2_io_V_wire_en_22[4'hd];
  assign T1102 = ArrayRowModule_2_io_V_wire_en_22[4'he];
  assign T1103 = ArrayRowModule_2_io_V_wire_en_22[4'hf];
  assign T1104 = ArrayRowModule_3_io_V_wire_en_0[1'h0];
  assign T1105 = ArrayRowModule_3_io_V_wire_en_0[1'h1];
  assign T1106 = ArrayRowModule_3_io_V_wire_en_0[2'h2];
  assign T1107 = ArrayRowModule_3_io_V_wire_en_0[2'h3];
  assign T1108 = ArrayRowModule_3_io_V_wire_en_0[3'h4];
  assign T1109 = ArrayRowModule_3_io_V_wire_en_0[3'h5];
  assign T1110 = ArrayRowModule_3_io_V_wire_en_0[3'h6];
  assign T1111 = ArrayRowModule_3_io_V_wire_en_0[3'h7];
  assign T1112 = ArrayRowModule_3_io_V_wire_en_0[4'h8];
  assign T1113 = ArrayRowModule_3_io_V_wire_en_0[4'h9];
  assign T1114 = ArrayRowModule_3_io_V_wire_en_0[4'ha];
  assign T1115 = ArrayRowModule_3_io_V_wire_en_0[4'hb];
  assign T1116 = ArrayRowModule_3_io_V_wire_en_0[4'hc];
  assign T1117 = ArrayRowModule_3_io_V_wire_en_0[4'hd];
  assign T1118 = ArrayRowModule_3_io_V_wire_en_0[4'he];
  assign T1119 = ArrayRowModule_3_io_V_wire_en_0[4'hf];
  assign T1120 = ArrayRowModule_3_io_V_wire_en_1[1'h0];
  assign T1121 = ArrayRowModule_3_io_V_wire_en_1[1'h1];
  assign T1122 = ArrayRowModule_3_io_V_wire_en_1[2'h2];
  assign T1123 = ArrayRowModule_3_io_V_wire_en_1[2'h3];
  assign T1124 = ArrayRowModule_3_io_V_wire_en_1[3'h4];
  assign T1125 = ArrayRowModule_3_io_V_wire_en_1[3'h5];
  assign T1126 = ArrayRowModule_3_io_V_wire_en_1[3'h6];
  assign T1127 = ArrayRowModule_3_io_V_wire_en_1[3'h7];
  assign T1128 = ArrayRowModule_3_io_V_wire_en_1[4'h8];
  assign T1129 = ArrayRowModule_3_io_V_wire_en_1[4'h9];
  assign T1130 = ArrayRowModule_3_io_V_wire_en_1[4'ha];
  assign T1131 = ArrayRowModule_3_io_V_wire_en_1[4'hb];
  assign T1132 = ArrayRowModule_3_io_V_wire_en_1[4'hc];
  assign T1133 = ArrayRowModule_3_io_V_wire_en_1[4'hd];
  assign T1134 = ArrayRowModule_3_io_V_wire_en_1[4'he];
  assign T1135 = ArrayRowModule_3_io_V_wire_en_1[4'hf];
  assign T1136 = ArrayRowModule_3_io_V_wire_en_2[1'h0];
  assign T1137 = ArrayRowModule_3_io_V_wire_en_2[1'h1];
  assign T1138 = ArrayRowModule_3_io_V_wire_en_2[2'h2];
  assign T1139 = ArrayRowModule_3_io_V_wire_en_2[2'h3];
  assign T1140 = ArrayRowModule_3_io_V_wire_en_2[3'h4];
  assign T1141 = ArrayRowModule_3_io_V_wire_en_2[3'h5];
  assign T1142 = ArrayRowModule_3_io_V_wire_en_2[3'h6];
  assign T1143 = ArrayRowModule_3_io_V_wire_en_2[3'h7];
  assign T1144 = ArrayRowModule_3_io_V_wire_en_2[4'h8];
  assign T1145 = ArrayRowModule_3_io_V_wire_en_2[4'h9];
  assign T1146 = ArrayRowModule_3_io_V_wire_en_2[4'ha];
  assign T1147 = ArrayRowModule_3_io_V_wire_en_2[4'hb];
  assign T1148 = ArrayRowModule_3_io_V_wire_en_2[4'hc];
  assign T1149 = ArrayRowModule_3_io_V_wire_en_2[4'hd];
  assign T1150 = ArrayRowModule_3_io_V_wire_en_2[4'he];
  assign T1151 = ArrayRowModule_3_io_V_wire_en_2[4'hf];
  assign T1152 = ArrayRowModule_3_io_V_wire_en_3[1'h0];
  assign T1153 = ArrayRowModule_3_io_V_wire_en_3[1'h1];
  assign T1154 = ArrayRowModule_3_io_V_wire_en_3[2'h2];
  assign T1155 = ArrayRowModule_3_io_V_wire_en_3[2'h3];
  assign T1156 = ArrayRowModule_3_io_V_wire_en_3[3'h4];
  assign T1157 = ArrayRowModule_3_io_V_wire_en_3[3'h5];
  assign T1158 = ArrayRowModule_3_io_V_wire_en_3[3'h6];
  assign T1159 = ArrayRowModule_3_io_V_wire_en_3[3'h7];
  assign T1160 = ArrayRowModule_3_io_V_wire_en_3[4'h8];
  assign T1161 = ArrayRowModule_3_io_V_wire_en_3[4'h9];
  assign T1162 = ArrayRowModule_3_io_V_wire_en_3[4'ha];
  assign T1163 = ArrayRowModule_3_io_V_wire_en_3[4'hb];
  assign T1164 = ArrayRowModule_3_io_V_wire_en_3[4'hc];
  assign T1165 = ArrayRowModule_3_io_V_wire_en_3[4'hd];
  assign T1166 = ArrayRowModule_3_io_V_wire_en_3[4'he];
  assign T1167 = ArrayRowModule_3_io_V_wire_en_3[4'hf];
  assign T1168 = ArrayRowModule_3_io_V_wire_en_4[1'h0];
  assign T1169 = ArrayRowModule_3_io_V_wire_en_4[1'h1];
  assign T1170 = ArrayRowModule_3_io_V_wire_en_4[2'h2];
  assign T1171 = ArrayRowModule_3_io_V_wire_en_4[2'h3];
  assign T1172 = ArrayRowModule_3_io_V_wire_en_4[3'h4];
  assign T1173 = ArrayRowModule_3_io_V_wire_en_4[3'h5];
  assign T1174 = ArrayRowModule_3_io_V_wire_en_4[3'h6];
  assign T1175 = ArrayRowModule_3_io_V_wire_en_4[3'h7];
  assign T1176 = ArrayRowModule_3_io_V_wire_en_4[4'h8];
  assign T1177 = ArrayRowModule_3_io_V_wire_en_4[4'h9];
  assign T1178 = ArrayRowModule_3_io_V_wire_en_4[4'ha];
  assign T1179 = ArrayRowModule_3_io_V_wire_en_4[4'hb];
  assign T1180 = ArrayRowModule_3_io_V_wire_en_4[4'hc];
  assign T1181 = ArrayRowModule_3_io_V_wire_en_4[4'hd];
  assign T1182 = ArrayRowModule_3_io_V_wire_en_4[4'he];
  assign T1183 = ArrayRowModule_3_io_V_wire_en_4[4'hf];
  assign T1184 = ArrayRowModule_3_io_V_wire_en_5[1'h0];
  assign T1185 = ArrayRowModule_3_io_V_wire_en_5[1'h1];
  assign T1186 = ArrayRowModule_3_io_V_wire_en_5[2'h2];
  assign T1187 = ArrayRowModule_3_io_V_wire_en_5[2'h3];
  assign T1188 = ArrayRowModule_3_io_V_wire_en_5[3'h4];
  assign T1189 = ArrayRowModule_3_io_V_wire_en_5[3'h5];
  assign T1190 = ArrayRowModule_3_io_V_wire_en_5[3'h6];
  assign T1191 = ArrayRowModule_3_io_V_wire_en_5[3'h7];
  assign T1192 = ArrayRowModule_3_io_V_wire_en_5[4'h8];
  assign T1193 = ArrayRowModule_3_io_V_wire_en_5[4'h9];
  assign T1194 = ArrayRowModule_3_io_V_wire_en_5[4'ha];
  assign T1195 = ArrayRowModule_3_io_V_wire_en_5[4'hb];
  assign T1196 = ArrayRowModule_3_io_V_wire_en_5[4'hc];
  assign T1197 = ArrayRowModule_3_io_V_wire_en_5[4'hd];
  assign T1198 = ArrayRowModule_3_io_V_wire_en_5[4'he];
  assign T1199 = ArrayRowModule_3_io_V_wire_en_5[4'hf];
  assign T1200 = ArrayRowModule_3_io_V_wire_en_6[1'h0];
  assign T1201 = ArrayRowModule_3_io_V_wire_en_6[1'h1];
  assign T1202 = ArrayRowModule_3_io_V_wire_en_6[2'h2];
  assign T1203 = ArrayRowModule_3_io_V_wire_en_6[2'h3];
  assign T1204 = ArrayRowModule_3_io_V_wire_en_6[3'h4];
  assign T1205 = ArrayRowModule_3_io_V_wire_en_6[3'h5];
  assign T1206 = ArrayRowModule_3_io_V_wire_en_6[3'h6];
  assign T1207 = ArrayRowModule_3_io_V_wire_en_6[3'h7];
  assign T1208 = ArrayRowModule_3_io_V_wire_en_6[4'h8];
  assign T1209 = ArrayRowModule_3_io_V_wire_en_6[4'h9];
  assign T1210 = ArrayRowModule_3_io_V_wire_en_6[4'ha];
  assign T1211 = ArrayRowModule_3_io_V_wire_en_6[4'hb];
  assign T1212 = ArrayRowModule_3_io_V_wire_en_6[4'hc];
  assign T1213 = ArrayRowModule_3_io_V_wire_en_6[4'hd];
  assign T1214 = ArrayRowModule_3_io_V_wire_en_6[4'he];
  assign T1215 = ArrayRowModule_3_io_V_wire_en_6[4'hf];
  assign T1216 = ArrayRowModule_3_io_V_wire_en_7[1'h0];
  assign T1217 = ArrayRowModule_3_io_V_wire_en_7[1'h1];
  assign T1218 = ArrayRowModule_3_io_V_wire_en_7[2'h2];
  assign T1219 = ArrayRowModule_3_io_V_wire_en_7[2'h3];
  assign T1220 = ArrayRowModule_3_io_V_wire_en_7[3'h4];
  assign T1221 = ArrayRowModule_3_io_V_wire_en_7[3'h5];
  assign T1222 = ArrayRowModule_3_io_V_wire_en_7[3'h6];
  assign T1223 = ArrayRowModule_3_io_V_wire_en_7[3'h7];
  assign T1224 = ArrayRowModule_3_io_V_wire_en_7[4'h8];
  assign T1225 = ArrayRowModule_3_io_V_wire_en_7[4'h9];
  assign T1226 = ArrayRowModule_3_io_V_wire_en_7[4'ha];
  assign T1227 = ArrayRowModule_3_io_V_wire_en_7[4'hb];
  assign T1228 = ArrayRowModule_3_io_V_wire_en_7[4'hc];
  assign T1229 = ArrayRowModule_3_io_V_wire_en_7[4'hd];
  assign T1230 = ArrayRowModule_3_io_V_wire_en_7[4'he];
  assign T1231 = ArrayRowModule_3_io_V_wire_en_7[4'hf];
  assign T1232 = ArrayRowModule_3_io_V_wire_en_8[1'h0];
  assign T1233 = ArrayRowModule_3_io_V_wire_en_8[1'h1];
  assign T1234 = ArrayRowModule_3_io_V_wire_en_8[2'h2];
  assign T1235 = ArrayRowModule_3_io_V_wire_en_8[2'h3];
  assign T1236 = ArrayRowModule_3_io_V_wire_en_8[3'h4];
  assign T1237 = ArrayRowModule_3_io_V_wire_en_8[3'h5];
  assign T1238 = ArrayRowModule_3_io_V_wire_en_8[3'h6];
  assign T1239 = ArrayRowModule_3_io_V_wire_en_8[3'h7];
  assign T1240 = ArrayRowModule_3_io_V_wire_en_8[4'h8];
  assign T1241 = ArrayRowModule_3_io_V_wire_en_8[4'h9];
  assign T1242 = ArrayRowModule_3_io_V_wire_en_8[4'ha];
  assign T1243 = ArrayRowModule_3_io_V_wire_en_8[4'hb];
  assign T1244 = ArrayRowModule_3_io_V_wire_en_8[4'hc];
  assign T1245 = ArrayRowModule_3_io_V_wire_en_8[4'hd];
  assign T1246 = ArrayRowModule_3_io_V_wire_en_8[4'he];
  assign T1247 = ArrayRowModule_3_io_V_wire_en_8[4'hf];
  assign T1248 = ArrayRowModule_3_io_V_wire_en_9[1'h0];
  assign T1249 = ArrayRowModule_3_io_V_wire_en_9[1'h1];
  assign T1250 = ArrayRowModule_3_io_V_wire_en_9[2'h2];
  assign T1251 = ArrayRowModule_3_io_V_wire_en_9[2'h3];
  assign T1252 = ArrayRowModule_3_io_V_wire_en_9[3'h4];
  assign T1253 = ArrayRowModule_3_io_V_wire_en_9[3'h5];
  assign T1254 = ArrayRowModule_3_io_V_wire_en_9[3'h6];
  assign T1255 = ArrayRowModule_3_io_V_wire_en_9[3'h7];
  assign T1256 = ArrayRowModule_3_io_V_wire_en_9[4'h8];
  assign T1257 = ArrayRowModule_3_io_V_wire_en_9[4'h9];
  assign T1258 = ArrayRowModule_3_io_V_wire_en_9[4'ha];
  assign T1259 = ArrayRowModule_3_io_V_wire_en_9[4'hb];
  assign T1260 = ArrayRowModule_3_io_V_wire_en_9[4'hc];
  assign T1261 = ArrayRowModule_3_io_V_wire_en_9[4'hd];
  assign T1262 = ArrayRowModule_3_io_V_wire_en_9[4'he];
  assign T1263 = ArrayRowModule_3_io_V_wire_en_9[4'hf];
  assign T1264 = ArrayRowModule_3_io_V_wire_en_10[1'h0];
  assign T1265 = ArrayRowModule_3_io_V_wire_en_10[1'h1];
  assign T1266 = ArrayRowModule_3_io_V_wire_en_10[2'h2];
  assign T1267 = ArrayRowModule_3_io_V_wire_en_10[2'h3];
  assign T1268 = ArrayRowModule_3_io_V_wire_en_10[3'h4];
  assign T1269 = ArrayRowModule_3_io_V_wire_en_10[3'h5];
  assign T1270 = ArrayRowModule_3_io_V_wire_en_10[3'h6];
  assign T1271 = ArrayRowModule_3_io_V_wire_en_10[3'h7];
  assign T1272 = ArrayRowModule_3_io_V_wire_en_10[4'h8];
  assign T1273 = ArrayRowModule_3_io_V_wire_en_10[4'h9];
  assign T1274 = ArrayRowModule_3_io_V_wire_en_10[4'ha];
  assign T1275 = ArrayRowModule_3_io_V_wire_en_10[4'hb];
  assign T1276 = ArrayRowModule_3_io_V_wire_en_10[4'hc];
  assign T1277 = ArrayRowModule_3_io_V_wire_en_10[4'hd];
  assign T1278 = ArrayRowModule_3_io_V_wire_en_10[4'he];
  assign T1279 = ArrayRowModule_3_io_V_wire_en_10[4'hf];
  assign T1280 = ArrayRowModule_3_io_V_wire_en_11[1'h0];
  assign T1281 = ArrayRowModule_3_io_V_wire_en_11[1'h1];
  assign T1282 = ArrayRowModule_3_io_V_wire_en_11[2'h2];
  assign T1283 = ArrayRowModule_3_io_V_wire_en_11[2'h3];
  assign T1284 = ArrayRowModule_3_io_V_wire_en_11[3'h4];
  assign T1285 = ArrayRowModule_3_io_V_wire_en_11[3'h5];
  assign T1286 = ArrayRowModule_3_io_V_wire_en_11[3'h6];
  assign T1287 = ArrayRowModule_3_io_V_wire_en_11[3'h7];
  assign T1288 = ArrayRowModule_3_io_V_wire_en_11[4'h8];
  assign T1289 = ArrayRowModule_3_io_V_wire_en_11[4'h9];
  assign T1290 = ArrayRowModule_3_io_V_wire_en_11[4'ha];
  assign T1291 = ArrayRowModule_3_io_V_wire_en_11[4'hb];
  assign T1292 = ArrayRowModule_3_io_V_wire_en_11[4'hc];
  assign T1293 = ArrayRowModule_3_io_V_wire_en_11[4'hd];
  assign T1294 = ArrayRowModule_3_io_V_wire_en_11[4'he];
  assign T1295 = ArrayRowModule_3_io_V_wire_en_11[4'hf];
  assign T1296 = ArrayRowModule_3_io_V_wire_en_12[1'h0];
  assign T1297 = ArrayRowModule_3_io_V_wire_en_12[1'h1];
  assign T1298 = ArrayRowModule_3_io_V_wire_en_12[2'h2];
  assign T1299 = ArrayRowModule_3_io_V_wire_en_12[2'h3];
  assign T1300 = ArrayRowModule_3_io_V_wire_en_12[3'h4];
  assign T1301 = ArrayRowModule_3_io_V_wire_en_12[3'h5];
  assign T1302 = ArrayRowModule_3_io_V_wire_en_12[3'h6];
  assign T1303 = ArrayRowModule_3_io_V_wire_en_12[3'h7];
  assign T1304 = ArrayRowModule_3_io_V_wire_en_12[4'h8];
  assign T1305 = ArrayRowModule_3_io_V_wire_en_12[4'h9];
  assign T1306 = ArrayRowModule_3_io_V_wire_en_12[4'ha];
  assign T1307 = ArrayRowModule_3_io_V_wire_en_12[4'hb];
  assign T1308 = ArrayRowModule_3_io_V_wire_en_12[4'hc];
  assign T1309 = ArrayRowModule_3_io_V_wire_en_12[4'hd];
  assign T1310 = ArrayRowModule_3_io_V_wire_en_12[4'he];
  assign T1311 = ArrayRowModule_3_io_V_wire_en_12[4'hf];
  assign T1312 = ArrayRowModule_3_io_V_wire_en_13[1'h0];
  assign T1313 = ArrayRowModule_3_io_V_wire_en_13[1'h1];
  assign T1314 = ArrayRowModule_3_io_V_wire_en_13[2'h2];
  assign T1315 = ArrayRowModule_3_io_V_wire_en_13[2'h3];
  assign T1316 = ArrayRowModule_3_io_V_wire_en_13[3'h4];
  assign T1317 = ArrayRowModule_3_io_V_wire_en_13[3'h5];
  assign T1318 = ArrayRowModule_3_io_V_wire_en_13[3'h6];
  assign T1319 = ArrayRowModule_3_io_V_wire_en_13[3'h7];
  assign T1320 = ArrayRowModule_3_io_V_wire_en_13[4'h8];
  assign T1321 = ArrayRowModule_3_io_V_wire_en_13[4'h9];
  assign T1322 = ArrayRowModule_3_io_V_wire_en_13[4'ha];
  assign T1323 = ArrayRowModule_3_io_V_wire_en_13[4'hb];
  assign T1324 = ArrayRowModule_3_io_V_wire_en_13[4'hc];
  assign T1325 = ArrayRowModule_3_io_V_wire_en_13[4'hd];
  assign T1326 = ArrayRowModule_3_io_V_wire_en_13[4'he];
  assign T1327 = ArrayRowModule_3_io_V_wire_en_13[4'hf];
  assign T1328 = ArrayRowModule_3_io_V_wire_en_14[1'h0];
  assign T1329 = ArrayRowModule_3_io_V_wire_en_14[1'h1];
  assign T1330 = ArrayRowModule_3_io_V_wire_en_14[2'h2];
  assign T1331 = ArrayRowModule_3_io_V_wire_en_14[2'h3];
  assign T1332 = ArrayRowModule_3_io_V_wire_en_14[3'h4];
  assign T1333 = ArrayRowModule_3_io_V_wire_en_14[3'h5];
  assign T1334 = ArrayRowModule_3_io_V_wire_en_14[3'h6];
  assign T1335 = ArrayRowModule_3_io_V_wire_en_14[3'h7];
  assign T1336 = ArrayRowModule_3_io_V_wire_en_14[4'h8];
  assign T1337 = ArrayRowModule_3_io_V_wire_en_14[4'h9];
  assign T1338 = ArrayRowModule_3_io_V_wire_en_14[4'ha];
  assign T1339 = ArrayRowModule_3_io_V_wire_en_14[4'hb];
  assign T1340 = ArrayRowModule_3_io_V_wire_en_14[4'hc];
  assign T1341 = ArrayRowModule_3_io_V_wire_en_14[4'hd];
  assign T1342 = ArrayRowModule_3_io_V_wire_en_14[4'he];
  assign T1343 = ArrayRowModule_3_io_V_wire_en_14[4'hf];
  assign T1344 = ArrayRowModule_3_io_V_wire_en_15[1'h0];
  assign T1345 = ArrayRowModule_3_io_V_wire_en_15[1'h1];
  assign T1346 = ArrayRowModule_3_io_V_wire_en_15[2'h2];
  assign T1347 = ArrayRowModule_3_io_V_wire_en_15[2'h3];
  assign T1348 = ArrayRowModule_3_io_V_wire_en_15[3'h4];
  assign T1349 = ArrayRowModule_3_io_V_wire_en_15[3'h5];
  assign T1350 = ArrayRowModule_3_io_V_wire_en_15[3'h6];
  assign T1351 = ArrayRowModule_3_io_V_wire_en_15[3'h7];
  assign T1352 = ArrayRowModule_3_io_V_wire_en_15[4'h8];
  assign T1353 = ArrayRowModule_3_io_V_wire_en_15[4'h9];
  assign T1354 = ArrayRowModule_3_io_V_wire_en_15[4'ha];
  assign T1355 = ArrayRowModule_3_io_V_wire_en_15[4'hb];
  assign T1356 = ArrayRowModule_3_io_V_wire_en_15[4'hc];
  assign T1357 = ArrayRowModule_3_io_V_wire_en_15[4'hd];
  assign T1358 = ArrayRowModule_3_io_V_wire_en_15[4'he];
  assign T1359 = ArrayRowModule_3_io_V_wire_en_15[4'hf];
  assign T1360 = ArrayRowModule_3_io_V_wire_en_16[1'h0];
  assign T1361 = ArrayRowModule_3_io_V_wire_en_16[1'h1];
  assign T1362 = ArrayRowModule_3_io_V_wire_en_16[2'h2];
  assign T1363 = ArrayRowModule_3_io_V_wire_en_16[2'h3];
  assign T1364 = ArrayRowModule_3_io_V_wire_en_16[3'h4];
  assign T1365 = ArrayRowModule_3_io_V_wire_en_16[3'h5];
  assign T1366 = ArrayRowModule_3_io_V_wire_en_16[3'h6];
  assign T1367 = ArrayRowModule_3_io_V_wire_en_16[3'h7];
  assign T1368 = ArrayRowModule_3_io_V_wire_en_16[4'h8];
  assign T1369 = ArrayRowModule_3_io_V_wire_en_16[4'h9];
  assign T1370 = ArrayRowModule_3_io_V_wire_en_16[4'ha];
  assign T1371 = ArrayRowModule_3_io_V_wire_en_16[4'hb];
  assign T1372 = ArrayRowModule_3_io_V_wire_en_16[4'hc];
  assign T1373 = ArrayRowModule_3_io_V_wire_en_16[4'hd];
  assign T1374 = ArrayRowModule_3_io_V_wire_en_16[4'he];
  assign T1375 = ArrayRowModule_3_io_V_wire_en_16[4'hf];
  assign T1376 = ArrayRowModule_3_io_V_wire_en_17[1'h0];
  assign T1377 = ArrayRowModule_3_io_V_wire_en_17[1'h1];
  assign T1378 = ArrayRowModule_3_io_V_wire_en_17[2'h2];
  assign T1379 = ArrayRowModule_3_io_V_wire_en_17[2'h3];
  assign T1380 = ArrayRowModule_3_io_V_wire_en_17[3'h4];
  assign T1381 = ArrayRowModule_3_io_V_wire_en_17[3'h5];
  assign T1382 = ArrayRowModule_3_io_V_wire_en_17[3'h6];
  assign T1383 = ArrayRowModule_3_io_V_wire_en_17[3'h7];
  assign T1384 = ArrayRowModule_3_io_V_wire_en_17[4'h8];
  assign T1385 = ArrayRowModule_3_io_V_wire_en_17[4'h9];
  assign T1386 = ArrayRowModule_3_io_V_wire_en_17[4'ha];
  assign T1387 = ArrayRowModule_3_io_V_wire_en_17[4'hb];
  assign T1388 = ArrayRowModule_3_io_V_wire_en_17[4'hc];
  assign T1389 = ArrayRowModule_3_io_V_wire_en_17[4'hd];
  assign T1390 = ArrayRowModule_3_io_V_wire_en_17[4'he];
  assign T1391 = ArrayRowModule_3_io_V_wire_en_17[4'hf];
  assign T1392 = ArrayRowModule_3_io_V_wire_en_18[1'h0];
  assign T1393 = ArrayRowModule_3_io_V_wire_en_18[1'h1];
  assign T1394 = ArrayRowModule_3_io_V_wire_en_18[2'h2];
  assign T1395 = ArrayRowModule_3_io_V_wire_en_18[2'h3];
  assign T1396 = ArrayRowModule_3_io_V_wire_en_18[3'h4];
  assign T1397 = ArrayRowModule_3_io_V_wire_en_18[3'h5];
  assign T1398 = ArrayRowModule_3_io_V_wire_en_18[3'h6];
  assign T1399 = ArrayRowModule_3_io_V_wire_en_18[3'h7];
  assign T1400 = ArrayRowModule_3_io_V_wire_en_18[4'h8];
  assign T1401 = ArrayRowModule_3_io_V_wire_en_18[4'h9];
  assign T1402 = ArrayRowModule_3_io_V_wire_en_18[4'ha];
  assign T1403 = ArrayRowModule_3_io_V_wire_en_18[4'hb];
  assign T1404 = ArrayRowModule_3_io_V_wire_en_18[4'hc];
  assign T1405 = ArrayRowModule_3_io_V_wire_en_18[4'hd];
  assign T1406 = ArrayRowModule_3_io_V_wire_en_18[4'he];
  assign T1407 = ArrayRowModule_3_io_V_wire_en_18[4'hf];
  assign T1408 = ArrayRowModule_3_io_V_wire_en_19[1'h0];
  assign T1409 = ArrayRowModule_3_io_V_wire_en_19[1'h1];
  assign T1410 = ArrayRowModule_3_io_V_wire_en_19[2'h2];
  assign T1411 = ArrayRowModule_3_io_V_wire_en_19[2'h3];
  assign T1412 = ArrayRowModule_3_io_V_wire_en_19[3'h4];
  assign T1413 = ArrayRowModule_3_io_V_wire_en_19[3'h5];
  assign T1414 = ArrayRowModule_3_io_V_wire_en_19[3'h6];
  assign T1415 = ArrayRowModule_3_io_V_wire_en_19[3'h7];
  assign T1416 = ArrayRowModule_3_io_V_wire_en_19[4'h8];
  assign T1417 = ArrayRowModule_3_io_V_wire_en_19[4'h9];
  assign T1418 = ArrayRowModule_3_io_V_wire_en_19[4'ha];
  assign T1419 = ArrayRowModule_3_io_V_wire_en_19[4'hb];
  assign T1420 = ArrayRowModule_3_io_V_wire_en_19[4'hc];
  assign T1421 = ArrayRowModule_3_io_V_wire_en_19[4'hd];
  assign T1422 = ArrayRowModule_3_io_V_wire_en_19[4'he];
  assign T1423 = ArrayRowModule_3_io_V_wire_en_19[4'hf];
  assign T1424 = ArrayRowModule_3_io_V_wire_en_20[1'h0];
  assign T1425 = ArrayRowModule_3_io_V_wire_en_20[1'h1];
  assign T1426 = ArrayRowModule_3_io_V_wire_en_20[2'h2];
  assign T1427 = ArrayRowModule_3_io_V_wire_en_20[2'h3];
  assign T1428 = ArrayRowModule_3_io_V_wire_en_20[3'h4];
  assign T1429 = ArrayRowModule_3_io_V_wire_en_20[3'h5];
  assign T1430 = ArrayRowModule_3_io_V_wire_en_20[3'h6];
  assign T1431 = ArrayRowModule_3_io_V_wire_en_20[3'h7];
  assign T1432 = ArrayRowModule_3_io_V_wire_en_20[4'h8];
  assign T1433 = ArrayRowModule_3_io_V_wire_en_20[4'h9];
  assign T1434 = ArrayRowModule_3_io_V_wire_en_20[4'ha];
  assign T1435 = ArrayRowModule_3_io_V_wire_en_20[4'hb];
  assign T1436 = ArrayRowModule_3_io_V_wire_en_20[4'hc];
  assign T1437 = ArrayRowModule_3_io_V_wire_en_20[4'hd];
  assign T1438 = ArrayRowModule_3_io_V_wire_en_20[4'he];
  assign T1439 = ArrayRowModule_3_io_V_wire_en_20[4'hf];
  assign T1440 = ArrayRowModule_3_io_V_wire_en_21[1'h0];
  assign T1441 = ArrayRowModule_3_io_V_wire_en_21[1'h1];
  assign T1442 = ArrayRowModule_3_io_V_wire_en_21[2'h2];
  assign T1443 = ArrayRowModule_3_io_V_wire_en_21[2'h3];
  assign T1444 = ArrayRowModule_3_io_V_wire_en_21[3'h4];
  assign T1445 = ArrayRowModule_3_io_V_wire_en_21[3'h5];
  assign T1446 = ArrayRowModule_3_io_V_wire_en_21[3'h6];
  assign T1447 = ArrayRowModule_3_io_V_wire_en_21[3'h7];
  assign T1448 = ArrayRowModule_3_io_V_wire_en_21[4'h8];
  assign T1449 = ArrayRowModule_3_io_V_wire_en_21[4'h9];
  assign T1450 = ArrayRowModule_3_io_V_wire_en_21[4'ha];
  assign T1451 = ArrayRowModule_3_io_V_wire_en_21[4'hb];
  assign T1452 = ArrayRowModule_3_io_V_wire_en_21[4'hc];
  assign T1453 = ArrayRowModule_3_io_V_wire_en_21[4'hd];
  assign T1454 = ArrayRowModule_3_io_V_wire_en_21[4'he];
  assign T1455 = ArrayRowModule_3_io_V_wire_en_21[4'hf];
  assign T1456 = ArrayRowModule_3_io_V_wire_en_22[1'h0];
  assign T1457 = ArrayRowModule_3_io_V_wire_en_22[1'h1];
  assign T1458 = ArrayRowModule_3_io_V_wire_en_22[2'h2];
  assign T1459 = ArrayRowModule_3_io_V_wire_en_22[2'h3];
  assign T1460 = ArrayRowModule_3_io_V_wire_en_22[3'h4];
  assign T1461 = ArrayRowModule_3_io_V_wire_en_22[3'h5];
  assign T1462 = ArrayRowModule_3_io_V_wire_en_22[3'h6];
  assign T1463 = ArrayRowModule_3_io_V_wire_en_22[3'h7];
  assign T1464 = ArrayRowModule_3_io_V_wire_en_22[4'h8];
  assign T1465 = ArrayRowModule_3_io_V_wire_en_22[4'h9];
  assign T1466 = ArrayRowModule_3_io_V_wire_en_22[4'ha];
  assign T1467 = ArrayRowModule_3_io_V_wire_en_22[4'hb];
  assign T1468 = ArrayRowModule_3_io_V_wire_en_22[4'hc];
  assign T1469 = ArrayRowModule_3_io_V_wire_en_22[4'hd];
  assign T1470 = ArrayRowModule_3_io_V_wire_en_22[4'he];
  assign T1471 = ArrayRowModule_3_io_V_wire_en_22[4'hf];
  assign T1472 = row_en[2'h3];
  assign row_en = ConfigAddrDecoder_io_en;
  assign T1473 = row_en[2'h2];
  assign T1474 = row_en[1'h1];
  assign T1475 = row_en[1'h0];
  assign io_mem_bus_out_0 = ArrayRowModule_3_io_mem_bus_out_0;
  assign io_mem_bus_out_1 = ArrayRowModule_3_io_mem_bus_out_1;
  assign io_mem_bus_out_2 = ArrayRowModule_3_io_mem_bus_out_2;
  assign io_mem_bus_out_3 = ArrayRowModule_3_io_mem_bus_out_3;
  assign io_mem_bus_out_4 = ArrayRowModule_3_io_mem_bus_out_4;
  assign io_mem_bus_out_5 = ArrayRowModule_3_io_mem_bus_out_5;
  assign io_mem_bus_out_6 = ArrayRowModule_3_io_mem_bus_out_6;
  assign io_mem_bus_out_7 = ArrayRowModule_3_io_mem_bus_out_7;
  assign io_mem_bus_out_8 = ArrayRowModule_3_io_mem_bus_out_8;
  assign io_mem_bus_out_9 = ArrayRowModule_3_io_mem_bus_out_9;
  assign io_mem_bus_out_10 = ArrayRowModule_3_io_mem_bus_out_10;
  assign io_mem_bus_out_11 = ArrayRowModule_3_io_mem_bus_out_11;
  assign io_mem_bus_out_12 = ArrayRowModule_3_io_mem_bus_out_12;
  assign io_mem_bus_out_13 = ArrayRowModule_3_io_mem_bus_out_13;
  assign io_mem_bus_out_14 = ArrayRowModule_3_io_mem_bus_out_14;
  assign io_mem_bus_out_15 = ArrayRowModule_3_io_mem_bus_out_15;
  assign io_mem_bus_out_16 = ArrayRowModule_3_io_mem_bus_out_16;
  assign io_mem_bus_out_17 = ArrayRowModule_3_io_mem_bus_out_17;
  assign io_mem_bus_out_18 = ArrayRowModule_3_io_mem_bus_out_18;
  assign io_mem_bus_out_19 = ArrayRowModule_3_io_mem_bus_out_19;
  assign io_mem_bus_out_20 = ArrayRowModule_3_io_mem_bus_out_20;
  assign io_mem_bus_out_21 = ArrayRowModule_3_io_mem_bus_out_21;
  assign io_mem_bus_out_22 = ArrayRowModule_3_io_mem_bus_out_22;
  assign io_mem_bus_out_23 = ArrayRowModule_3_io_mem_bus_out_23;
  ConfigAddrDecoder ConfigAddrDecoder(
       .io_addr( io_addr ),
       .io_en( ConfigAddrDecoder_io_en )
  );
  ArrayRowModule ArrayRowModule(.clk(clk), .reset(reset),
       .io_V_wire_in_367( VwireModule_io_VwirePorts_0_22_15_out ),
       .io_V_wire_in_366( VwireModule_io_VwirePorts_0_22_14_out ),
       .io_V_wire_in_365( VwireModule_io_VwirePorts_0_22_13_out ),
       .io_V_wire_in_364( VwireModule_io_VwirePorts_0_22_12_out ),
       .io_V_wire_in_363( VwireModule_io_VwirePorts_0_22_11_out ),
       .io_V_wire_in_362( VwireModule_io_VwirePorts_0_22_10_out ),
       .io_V_wire_in_361( VwireModule_io_VwirePorts_0_22_9_out ),
       .io_V_wire_in_360( VwireModule_io_VwirePorts_0_22_8_out ),
       .io_V_wire_in_359( VwireModule_io_VwirePorts_0_22_7_out ),
       .io_V_wire_in_358( VwireModule_io_VwirePorts_0_22_6_out ),
       .io_V_wire_in_357( VwireModule_io_VwirePorts_0_22_5_out ),
       .io_V_wire_in_356( VwireModule_io_VwirePorts_0_22_4_out ),
       .io_V_wire_in_355( VwireModule_io_VwirePorts_0_22_3_out ),
       .io_V_wire_in_354( VwireModule_io_VwirePorts_0_22_2_out ),
       .io_V_wire_in_353( VwireModule_io_VwirePorts_0_22_1_out ),
       .io_V_wire_in_352( VwireModule_io_VwirePorts_0_22_0_out ),
       .io_V_wire_in_351( VwireModule_io_VwirePorts_0_21_15_out ),
       .io_V_wire_in_350( VwireModule_io_VwirePorts_0_21_14_out ),
       .io_V_wire_in_349( VwireModule_io_VwirePorts_0_21_13_out ),
       .io_V_wire_in_348( VwireModule_io_VwirePorts_0_21_12_out ),
       .io_V_wire_in_347( VwireModule_io_VwirePorts_0_21_11_out ),
       .io_V_wire_in_346( VwireModule_io_VwirePorts_0_21_10_out ),
       .io_V_wire_in_345( VwireModule_io_VwirePorts_0_21_9_out ),
       .io_V_wire_in_344( VwireModule_io_VwirePorts_0_21_8_out ),
       .io_V_wire_in_343( VwireModule_io_VwirePorts_0_21_7_out ),
       .io_V_wire_in_342( VwireModule_io_VwirePorts_0_21_6_out ),
       .io_V_wire_in_341( VwireModule_io_VwirePorts_0_21_5_out ),
       .io_V_wire_in_340( VwireModule_io_VwirePorts_0_21_4_out ),
       .io_V_wire_in_339( VwireModule_io_VwirePorts_0_21_3_out ),
       .io_V_wire_in_338( VwireModule_io_VwirePorts_0_21_2_out ),
       .io_V_wire_in_337( VwireModule_io_VwirePorts_0_21_1_out ),
       .io_V_wire_in_336( VwireModule_io_VwirePorts_0_21_0_out ),
       .io_V_wire_in_335( VwireModule_io_VwirePorts_0_20_15_out ),
       .io_V_wire_in_334( VwireModule_io_VwirePorts_0_20_14_out ),
       .io_V_wire_in_333( VwireModule_io_VwirePorts_0_20_13_out ),
       .io_V_wire_in_332( VwireModule_io_VwirePorts_0_20_12_out ),
       .io_V_wire_in_331( VwireModule_io_VwirePorts_0_20_11_out ),
       .io_V_wire_in_330( VwireModule_io_VwirePorts_0_20_10_out ),
       .io_V_wire_in_329( VwireModule_io_VwirePorts_0_20_9_out ),
       .io_V_wire_in_328( VwireModule_io_VwirePorts_0_20_8_out ),
       .io_V_wire_in_327( VwireModule_io_VwirePorts_0_20_7_out ),
       .io_V_wire_in_326( VwireModule_io_VwirePorts_0_20_6_out ),
       .io_V_wire_in_325( VwireModule_io_VwirePorts_0_20_5_out ),
       .io_V_wire_in_324( VwireModule_io_VwirePorts_0_20_4_out ),
       .io_V_wire_in_323( VwireModule_io_VwirePorts_0_20_3_out ),
       .io_V_wire_in_322( VwireModule_io_VwirePorts_0_20_2_out ),
       .io_V_wire_in_321( VwireModule_io_VwirePorts_0_20_1_out ),
       .io_V_wire_in_320( VwireModule_io_VwirePorts_0_20_0_out ),
       .io_V_wire_in_319( VwireModule_io_VwirePorts_0_19_15_out ),
       .io_V_wire_in_318( VwireModule_io_VwirePorts_0_19_14_out ),
       .io_V_wire_in_317( VwireModule_io_VwirePorts_0_19_13_out ),
       .io_V_wire_in_316( VwireModule_io_VwirePorts_0_19_12_out ),
       .io_V_wire_in_315( VwireModule_io_VwirePorts_0_19_11_out ),
       .io_V_wire_in_314( VwireModule_io_VwirePorts_0_19_10_out ),
       .io_V_wire_in_313( VwireModule_io_VwirePorts_0_19_9_out ),
       .io_V_wire_in_312( VwireModule_io_VwirePorts_0_19_8_out ),
       .io_V_wire_in_311( VwireModule_io_VwirePorts_0_19_7_out ),
       .io_V_wire_in_310( VwireModule_io_VwirePorts_0_19_6_out ),
       .io_V_wire_in_309( VwireModule_io_VwirePorts_0_19_5_out ),
       .io_V_wire_in_308( VwireModule_io_VwirePorts_0_19_4_out ),
       .io_V_wire_in_307( VwireModule_io_VwirePorts_0_19_3_out ),
       .io_V_wire_in_306( VwireModule_io_VwirePorts_0_19_2_out ),
       .io_V_wire_in_305( VwireModule_io_VwirePorts_0_19_1_out ),
       .io_V_wire_in_304( VwireModule_io_VwirePorts_0_19_0_out ),
       .io_V_wire_in_303( VwireModule_io_VwirePorts_0_18_15_out ),
       .io_V_wire_in_302( VwireModule_io_VwirePorts_0_18_14_out ),
       .io_V_wire_in_301( VwireModule_io_VwirePorts_0_18_13_out ),
       .io_V_wire_in_300( VwireModule_io_VwirePorts_0_18_12_out ),
       .io_V_wire_in_299( VwireModule_io_VwirePorts_0_18_11_out ),
       .io_V_wire_in_298( VwireModule_io_VwirePorts_0_18_10_out ),
       .io_V_wire_in_297( VwireModule_io_VwirePorts_0_18_9_out ),
       .io_V_wire_in_296( VwireModule_io_VwirePorts_0_18_8_out ),
       .io_V_wire_in_295( VwireModule_io_VwirePorts_0_18_7_out ),
       .io_V_wire_in_294( VwireModule_io_VwirePorts_0_18_6_out ),
       .io_V_wire_in_293( VwireModule_io_VwirePorts_0_18_5_out ),
       .io_V_wire_in_292( VwireModule_io_VwirePorts_0_18_4_out ),
       .io_V_wire_in_291( VwireModule_io_VwirePorts_0_18_3_out ),
       .io_V_wire_in_290( VwireModule_io_VwirePorts_0_18_2_out ),
       .io_V_wire_in_289( VwireModule_io_VwirePorts_0_18_1_out ),
       .io_V_wire_in_288( VwireModule_io_VwirePorts_0_18_0_out ),
       .io_V_wire_in_287( VwireModule_io_VwirePorts_0_17_15_out ),
       .io_V_wire_in_286( VwireModule_io_VwirePorts_0_17_14_out ),
       .io_V_wire_in_285( VwireModule_io_VwirePorts_0_17_13_out ),
       .io_V_wire_in_284( VwireModule_io_VwirePorts_0_17_12_out ),
       .io_V_wire_in_283( VwireModule_io_VwirePorts_0_17_11_out ),
       .io_V_wire_in_282( VwireModule_io_VwirePorts_0_17_10_out ),
       .io_V_wire_in_281( VwireModule_io_VwirePorts_0_17_9_out ),
       .io_V_wire_in_280( VwireModule_io_VwirePorts_0_17_8_out ),
       .io_V_wire_in_279( VwireModule_io_VwirePorts_0_17_7_out ),
       .io_V_wire_in_278( VwireModule_io_VwirePorts_0_17_6_out ),
       .io_V_wire_in_277( VwireModule_io_VwirePorts_0_17_5_out ),
       .io_V_wire_in_276( VwireModule_io_VwirePorts_0_17_4_out ),
       .io_V_wire_in_275( VwireModule_io_VwirePorts_0_17_3_out ),
       .io_V_wire_in_274( VwireModule_io_VwirePorts_0_17_2_out ),
       .io_V_wire_in_273( VwireModule_io_VwirePorts_0_17_1_out ),
       .io_V_wire_in_272( VwireModule_io_VwirePorts_0_17_0_out ),
       .io_V_wire_in_271( VwireModule_io_VwirePorts_0_16_15_out ),
       .io_V_wire_in_270( VwireModule_io_VwirePorts_0_16_14_out ),
       .io_V_wire_in_269( VwireModule_io_VwirePorts_0_16_13_out ),
       .io_V_wire_in_268( VwireModule_io_VwirePorts_0_16_12_out ),
       .io_V_wire_in_267( VwireModule_io_VwirePorts_0_16_11_out ),
       .io_V_wire_in_266( VwireModule_io_VwirePorts_0_16_10_out ),
       .io_V_wire_in_265( VwireModule_io_VwirePorts_0_16_9_out ),
       .io_V_wire_in_264( VwireModule_io_VwirePorts_0_16_8_out ),
       .io_V_wire_in_263( VwireModule_io_VwirePorts_0_16_7_out ),
       .io_V_wire_in_262( VwireModule_io_VwirePorts_0_16_6_out ),
       .io_V_wire_in_261( VwireModule_io_VwirePorts_0_16_5_out ),
       .io_V_wire_in_260( VwireModule_io_VwirePorts_0_16_4_out ),
       .io_V_wire_in_259( VwireModule_io_VwirePorts_0_16_3_out ),
       .io_V_wire_in_258( VwireModule_io_VwirePorts_0_16_2_out ),
       .io_V_wire_in_257( VwireModule_io_VwirePorts_0_16_1_out ),
       .io_V_wire_in_256( VwireModule_io_VwirePorts_0_16_0_out ),
       .io_V_wire_in_255( VwireModule_io_VwirePorts_0_15_15_out ),
       .io_V_wire_in_254( VwireModule_io_VwirePorts_0_15_14_out ),
       .io_V_wire_in_253( VwireModule_io_VwirePorts_0_15_13_out ),
       .io_V_wire_in_252( VwireModule_io_VwirePorts_0_15_12_out ),
       .io_V_wire_in_251( VwireModule_io_VwirePorts_0_15_11_out ),
       .io_V_wire_in_250( VwireModule_io_VwirePorts_0_15_10_out ),
       .io_V_wire_in_249( VwireModule_io_VwirePorts_0_15_9_out ),
       .io_V_wire_in_248( VwireModule_io_VwirePorts_0_15_8_out ),
       .io_V_wire_in_247( VwireModule_io_VwirePorts_0_15_7_out ),
       .io_V_wire_in_246( VwireModule_io_VwirePorts_0_15_6_out ),
       .io_V_wire_in_245( VwireModule_io_VwirePorts_0_15_5_out ),
       .io_V_wire_in_244( VwireModule_io_VwirePorts_0_15_4_out ),
       .io_V_wire_in_243( VwireModule_io_VwirePorts_0_15_3_out ),
       .io_V_wire_in_242( VwireModule_io_VwirePorts_0_15_2_out ),
       .io_V_wire_in_241( VwireModule_io_VwirePorts_0_15_1_out ),
       .io_V_wire_in_240( VwireModule_io_VwirePorts_0_15_0_out ),
       .io_V_wire_in_239( VwireModule_io_VwirePorts_0_14_15_out ),
       .io_V_wire_in_238( VwireModule_io_VwirePorts_0_14_14_out ),
       .io_V_wire_in_237( VwireModule_io_VwirePorts_0_14_13_out ),
       .io_V_wire_in_236( VwireModule_io_VwirePorts_0_14_12_out ),
       .io_V_wire_in_235( VwireModule_io_VwirePorts_0_14_11_out ),
       .io_V_wire_in_234( VwireModule_io_VwirePorts_0_14_10_out ),
       .io_V_wire_in_233( VwireModule_io_VwirePorts_0_14_9_out ),
       .io_V_wire_in_232( VwireModule_io_VwirePorts_0_14_8_out ),
       .io_V_wire_in_231( VwireModule_io_VwirePorts_0_14_7_out ),
       .io_V_wire_in_230( VwireModule_io_VwirePorts_0_14_6_out ),
       .io_V_wire_in_229( VwireModule_io_VwirePorts_0_14_5_out ),
       .io_V_wire_in_228( VwireModule_io_VwirePorts_0_14_4_out ),
       .io_V_wire_in_227( VwireModule_io_VwirePorts_0_14_3_out ),
       .io_V_wire_in_226( VwireModule_io_VwirePorts_0_14_2_out ),
       .io_V_wire_in_225( VwireModule_io_VwirePorts_0_14_1_out ),
       .io_V_wire_in_224( VwireModule_io_VwirePorts_0_14_0_out ),
       .io_V_wire_in_223( VwireModule_io_VwirePorts_0_13_15_out ),
       .io_V_wire_in_222( VwireModule_io_VwirePorts_0_13_14_out ),
       .io_V_wire_in_221( VwireModule_io_VwirePorts_0_13_13_out ),
       .io_V_wire_in_220( VwireModule_io_VwirePorts_0_13_12_out ),
       .io_V_wire_in_219( VwireModule_io_VwirePorts_0_13_11_out ),
       .io_V_wire_in_218( VwireModule_io_VwirePorts_0_13_10_out ),
       .io_V_wire_in_217( VwireModule_io_VwirePorts_0_13_9_out ),
       .io_V_wire_in_216( VwireModule_io_VwirePorts_0_13_8_out ),
       .io_V_wire_in_215( VwireModule_io_VwirePorts_0_13_7_out ),
       .io_V_wire_in_214( VwireModule_io_VwirePorts_0_13_6_out ),
       .io_V_wire_in_213( VwireModule_io_VwirePorts_0_13_5_out ),
       .io_V_wire_in_212( VwireModule_io_VwirePorts_0_13_4_out ),
       .io_V_wire_in_211( VwireModule_io_VwirePorts_0_13_3_out ),
       .io_V_wire_in_210( VwireModule_io_VwirePorts_0_13_2_out ),
       .io_V_wire_in_209( VwireModule_io_VwirePorts_0_13_1_out ),
       .io_V_wire_in_208( VwireModule_io_VwirePorts_0_13_0_out ),
       .io_V_wire_in_207( VwireModule_io_VwirePorts_0_12_15_out ),
       .io_V_wire_in_206( VwireModule_io_VwirePorts_0_12_14_out ),
       .io_V_wire_in_205( VwireModule_io_VwirePorts_0_12_13_out ),
       .io_V_wire_in_204( VwireModule_io_VwirePorts_0_12_12_out ),
       .io_V_wire_in_203( VwireModule_io_VwirePorts_0_12_11_out ),
       .io_V_wire_in_202( VwireModule_io_VwirePorts_0_12_10_out ),
       .io_V_wire_in_201( VwireModule_io_VwirePorts_0_12_9_out ),
       .io_V_wire_in_200( VwireModule_io_VwirePorts_0_12_8_out ),
       .io_V_wire_in_199( VwireModule_io_VwirePorts_0_12_7_out ),
       .io_V_wire_in_198( VwireModule_io_VwirePorts_0_12_6_out ),
       .io_V_wire_in_197( VwireModule_io_VwirePorts_0_12_5_out ),
       .io_V_wire_in_196( VwireModule_io_VwirePorts_0_12_4_out ),
       .io_V_wire_in_195( VwireModule_io_VwirePorts_0_12_3_out ),
       .io_V_wire_in_194( VwireModule_io_VwirePorts_0_12_2_out ),
       .io_V_wire_in_193( VwireModule_io_VwirePorts_0_12_1_out ),
       .io_V_wire_in_192( VwireModule_io_VwirePorts_0_12_0_out ),
       .io_V_wire_in_191( VwireModule_io_VwirePorts_0_11_15_out ),
       .io_V_wire_in_190( VwireModule_io_VwirePorts_0_11_14_out ),
       .io_V_wire_in_189( VwireModule_io_VwirePorts_0_11_13_out ),
       .io_V_wire_in_188( VwireModule_io_VwirePorts_0_11_12_out ),
       .io_V_wire_in_187( VwireModule_io_VwirePorts_0_11_11_out ),
       .io_V_wire_in_186( VwireModule_io_VwirePorts_0_11_10_out ),
       .io_V_wire_in_185( VwireModule_io_VwirePorts_0_11_9_out ),
       .io_V_wire_in_184( VwireModule_io_VwirePorts_0_11_8_out ),
       .io_V_wire_in_183( VwireModule_io_VwirePorts_0_11_7_out ),
       .io_V_wire_in_182( VwireModule_io_VwirePorts_0_11_6_out ),
       .io_V_wire_in_181( VwireModule_io_VwirePorts_0_11_5_out ),
       .io_V_wire_in_180( VwireModule_io_VwirePorts_0_11_4_out ),
       .io_V_wire_in_179( VwireModule_io_VwirePorts_0_11_3_out ),
       .io_V_wire_in_178( VwireModule_io_VwirePorts_0_11_2_out ),
       .io_V_wire_in_177( VwireModule_io_VwirePorts_0_11_1_out ),
       .io_V_wire_in_176( VwireModule_io_VwirePorts_0_11_0_out ),
       .io_V_wire_in_175( VwireModule_io_VwirePorts_0_10_15_out ),
       .io_V_wire_in_174( VwireModule_io_VwirePorts_0_10_14_out ),
       .io_V_wire_in_173( VwireModule_io_VwirePorts_0_10_13_out ),
       .io_V_wire_in_172( VwireModule_io_VwirePorts_0_10_12_out ),
       .io_V_wire_in_171( VwireModule_io_VwirePorts_0_10_11_out ),
       .io_V_wire_in_170( VwireModule_io_VwirePorts_0_10_10_out ),
       .io_V_wire_in_169( VwireModule_io_VwirePorts_0_10_9_out ),
       .io_V_wire_in_168( VwireModule_io_VwirePorts_0_10_8_out ),
       .io_V_wire_in_167( VwireModule_io_VwirePorts_0_10_7_out ),
       .io_V_wire_in_166( VwireModule_io_VwirePorts_0_10_6_out ),
       .io_V_wire_in_165( VwireModule_io_VwirePorts_0_10_5_out ),
       .io_V_wire_in_164( VwireModule_io_VwirePorts_0_10_4_out ),
       .io_V_wire_in_163( VwireModule_io_VwirePorts_0_10_3_out ),
       .io_V_wire_in_162( VwireModule_io_VwirePorts_0_10_2_out ),
       .io_V_wire_in_161( VwireModule_io_VwirePorts_0_10_1_out ),
       .io_V_wire_in_160( VwireModule_io_VwirePorts_0_10_0_out ),
       .io_V_wire_in_159( VwireModule_io_VwirePorts_0_9_15_out ),
       .io_V_wire_in_158( VwireModule_io_VwirePorts_0_9_14_out ),
       .io_V_wire_in_157( VwireModule_io_VwirePorts_0_9_13_out ),
       .io_V_wire_in_156( VwireModule_io_VwirePorts_0_9_12_out ),
       .io_V_wire_in_155( VwireModule_io_VwirePorts_0_9_11_out ),
       .io_V_wire_in_154( VwireModule_io_VwirePorts_0_9_10_out ),
       .io_V_wire_in_153( VwireModule_io_VwirePorts_0_9_9_out ),
       .io_V_wire_in_152( VwireModule_io_VwirePorts_0_9_8_out ),
       .io_V_wire_in_151( VwireModule_io_VwirePorts_0_9_7_out ),
       .io_V_wire_in_150( VwireModule_io_VwirePorts_0_9_6_out ),
       .io_V_wire_in_149( VwireModule_io_VwirePorts_0_9_5_out ),
       .io_V_wire_in_148( VwireModule_io_VwirePorts_0_9_4_out ),
       .io_V_wire_in_147( VwireModule_io_VwirePorts_0_9_3_out ),
       .io_V_wire_in_146( VwireModule_io_VwirePorts_0_9_2_out ),
       .io_V_wire_in_145( VwireModule_io_VwirePorts_0_9_1_out ),
       .io_V_wire_in_144( VwireModule_io_VwirePorts_0_9_0_out ),
       .io_V_wire_in_143( VwireModule_io_VwirePorts_0_8_15_out ),
       .io_V_wire_in_142( VwireModule_io_VwirePorts_0_8_14_out ),
       .io_V_wire_in_141( VwireModule_io_VwirePorts_0_8_13_out ),
       .io_V_wire_in_140( VwireModule_io_VwirePorts_0_8_12_out ),
       .io_V_wire_in_139( VwireModule_io_VwirePorts_0_8_11_out ),
       .io_V_wire_in_138( VwireModule_io_VwirePorts_0_8_10_out ),
       .io_V_wire_in_137( VwireModule_io_VwirePorts_0_8_9_out ),
       .io_V_wire_in_136( VwireModule_io_VwirePorts_0_8_8_out ),
       .io_V_wire_in_135( VwireModule_io_VwirePorts_0_8_7_out ),
       .io_V_wire_in_134( VwireModule_io_VwirePorts_0_8_6_out ),
       .io_V_wire_in_133( VwireModule_io_VwirePorts_0_8_5_out ),
       .io_V_wire_in_132( VwireModule_io_VwirePorts_0_8_4_out ),
       .io_V_wire_in_131( VwireModule_io_VwirePorts_0_8_3_out ),
       .io_V_wire_in_130( VwireModule_io_VwirePorts_0_8_2_out ),
       .io_V_wire_in_129( VwireModule_io_VwirePorts_0_8_1_out ),
       .io_V_wire_in_128( VwireModule_io_VwirePorts_0_8_0_out ),
       .io_V_wire_in_127( VwireModule_io_VwirePorts_0_7_15_out ),
       .io_V_wire_in_126( VwireModule_io_VwirePorts_0_7_14_out ),
       .io_V_wire_in_125( VwireModule_io_VwirePorts_0_7_13_out ),
       .io_V_wire_in_124( VwireModule_io_VwirePorts_0_7_12_out ),
       .io_V_wire_in_123( VwireModule_io_VwirePorts_0_7_11_out ),
       .io_V_wire_in_122( VwireModule_io_VwirePorts_0_7_10_out ),
       .io_V_wire_in_121( VwireModule_io_VwirePorts_0_7_9_out ),
       .io_V_wire_in_120( VwireModule_io_VwirePorts_0_7_8_out ),
       .io_V_wire_in_119( VwireModule_io_VwirePorts_0_7_7_out ),
       .io_V_wire_in_118( VwireModule_io_VwirePorts_0_7_6_out ),
       .io_V_wire_in_117( VwireModule_io_VwirePorts_0_7_5_out ),
       .io_V_wire_in_116( VwireModule_io_VwirePorts_0_7_4_out ),
       .io_V_wire_in_115( VwireModule_io_VwirePorts_0_7_3_out ),
       .io_V_wire_in_114( VwireModule_io_VwirePorts_0_7_2_out ),
       .io_V_wire_in_113( VwireModule_io_VwirePorts_0_7_1_out ),
       .io_V_wire_in_112( VwireModule_io_VwirePorts_0_7_0_out ),
       .io_V_wire_in_111( VwireModule_io_VwirePorts_0_6_15_out ),
       .io_V_wire_in_110( VwireModule_io_VwirePorts_0_6_14_out ),
       .io_V_wire_in_109( VwireModule_io_VwirePorts_0_6_13_out ),
       .io_V_wire_in_108( VwireModule_io_VwirePorts_0_6_12_out ),
       .io_V_wire_in_107( VwireModule_io_VwirePorts_0_6_11_out ),
       .io_V_wire_in_106( VwireModule_io_VwirePorts_0_6_10_out ),
       .io_V_wire_in_105( VwireModule_io_VwirePorts_0_6_9_out ),
       .io_V_wire_in_104( VwireModule_io_VwirePorts_0_6_8_out ),
       .io_V_wire_in_103( VwireModule_io_VwirePorts_0_6_7_out ),
       .io_V_wire_in_102( VwireModule_io_VwirePorts_0_6_6_out ),
       .io_V_wire_in_101( VwireModule_io_VwirePorts_0_6_5_out ),
       .io_V_wire_in_100( VwireModule_io_VwirePorts_0_6_4_out ),
       .io_V_wire_in_99( VwireModule_io_VwirePorts_0_6_3_out ),
       .io_V_wire_in_98( VwireModule_io_VwirePorts_0_6_2_out ),
       .io_V_wire_in_97( VwireModule_io_VwirePorts_0_6_1_out ),
       .io_V_wire_in_96( VwireModule_io_VwirePorts_0_6_0_out ),
       .io_V_wire_in_95( VwireModule_io_VwirePorts_0_5_15_out ),
       .io_V_wire_in_94( VwireModule_io_VwirePorts_0_5_14_out ),
       .io_V_wire_in_93( VwireModule_io_VwirePorts_0_5_13_out ),
       .io_V_wire_in_92( VwireModule_io_VwirePorts_0_5_12_out ),
       .io_V_wire_in_91( VwireModule_io_VwirePorts_0_5_11_out ),
       .io_V_wire_in_90( VwireModule_io_VwirePorts_0_5_10_out ),
       .io_V_wire_in_89( VwireModule_io_VwirePorts_0_5_9_out ),
       .io_V_wire_in_88( VwireModule_io_VwirePorts_0_5_8_out ),
       .io_V_wire_in_87( VwireModule_io_VwirePorts_0_5_7_out ),
       .io_V_wire_in_86( VwireModule_io_VwirePorts_0_5_6_out ),
       .io_V_wire_in_85( VwireModule_io_VwirePorts_0_5_5_out ),
       .io_V_wire_in_84( VwireModule_io_VwirePorts_0_5_4_out ),
       .io_V_wire_in_83( VwireModule_io_VwirePorts_0_5_3_out ),
       .io_V_wire_in_82( VwireModule_io_VwirePorts_0_5_2_out ),
       .io_V_wire_in_81( VwireModule_io_VwirePorts_0_5_1_out ),
       .io_V_wire_in_80( VwireModule_io_VwirePorts_0_5_0_out ),
       .io_V_wire_in_79( VwireModule_io_VwirePorts_0_4_15_out ),
       .io_V_wire_in_78( VwireModule_io_VwirePorts_0_4_14_out ),
       .io_V_wire_in_77( VwireModule_io_VwirePorts_0_4_13_out ),
       .io_V_wire_in_76( VwireModule_io_VwirePorts_0_4_12_out ),
       .io_V_wire_in_75( VwireModule_io_VwirePorts_0_4_11_out ),
       .io_V_wire_in_74( VwireModule_io_VwirePorts_0_4_10_out ),
       .io_V_wire_in_73( VwireModule_io_VwirePorts_0_4_9_out ),
       .io_V_wire_in_72( VwireModule_io_VwirePorts_0_4_8_out ),
       .io_V_wire_in_71( VwireModule_io_VwirePorts_0_4_7_out ),
       .io_V_wire_in_70( VwireModule_io_VwirePorts_0_4_6_out ),
       .io_V_wire_in_69( VwireModule_io_VwirePorts_0_4_5_out ),
       .io_V_wire_in_68( VwireModule_io_VwirePorts_0_4_4_out ),
       .io_V_wire_in_67( VwireModule_io_VwirePorts_0_4_3_out ),
       .io_V_wire_in_66( VwireModule_io_VwirePorts_0_4_2_out ),
       .io_V_wire_in_65( VwireModule_io_VwirePorts_0_4_1_out ),
       .io_V_wire_in_64( VwireModule_io_VwirePorts_0_4_0_out ),
       .io_V_wire_in_63( VwireModule_io_VwirePorts_0_3_15_out ),
       .io_V_wire_in_62( VwireModule_io_VwirePorts_0_3_14_out ),
       .io_V_wire_in_61( VwireModule_io_VwirePorts_0_3_13_out ),
       .io_V_wire_in_60( VwireModule_io_VwirePorts_0_3_12_out ),
       .io_V_wire_in_59( VwireModule_io_VwirePorts_0_3_11_out ),
       .io_V_wire_in_58( VwireModule_io_VwirePorts_0_3_10_out ),
       .io_V_wire_in_57( VwireModule_io_VwirePorts_0_3_9_out ),
       .io_V_wire_in_56( VwireModule_io_VwirePorts_0_3_8_out ),
       .io_V_wire_in_55( VwireModule_io_VwirePorts_0_3_7_out ),
       .io_V_wire_in_54( VwireModule_io_VwirePorts_0_3_6_out ),
       .io_V_wire_in_53( VwireModule_io_VwirePorts_0_3_5_out ),
       .io_V_wire_in_52( VwireModule_io_VwirePorts_0_3_4_out ),
       .io_V_wire_in_51( VwireModule_io_VwirePorts_0_3_3_out ),
       .io_V_wire_in_50( VwireModule_io_VwirePorts_0_3_2_out ),
       .io_V_wire_in_49( VwireModule_io_VwirePorts_0_3_1_out ),
       .io_V_wire_in_48( VwireModule_io_VwirePorts_0_3_0_out ),
       .io_V_wire_in_47( VwireModule_io_VwirePorts_0_2_15_out ),
       .io_V_wire_in_46( VwireModule_io_VwirePorts_0_2_14_out ),
       .io_V_wire_in_45( VwireModule_io_VwirePorts_0_2_13_out ),
       .io_V_wire_in_44( VwireModule_io_VwirePorts_0_2_12_out ),
       .io_V_wire_in_43( VwireModule_io_VwirePorts_0_2_11_out ),
       .io_V_wire_in_42( VwireModule_io_VwirePorts_0_2_10_out ),
       .io_V_wire_in_41( VwireModule_io_VwirePorts_0_2_9_out ),
       .io_V_wire_in_40( VwireModule_io_VwirePorts_0_2_8_out ),
       .io_V_wire_in_39( VwireModule_io_VwirePorts_0_2_7_out ),
       .io_V_wire_in_38( VwireModule_io_VwirePorts_0_2_6_out ),
       .io_V_wire_in_37( VwireModule_io_VwirePorts_0_2_5_out ),
       .io_V_wire_in_36( VwireModule_io_VwirePorts_0_2_4_out ),
       .io_V_wire_in_35( VwireModule_io_VwirePorts_0_2_3_out ),
       .io_V_wire_in_34( VwireModule_io_VwirePorts_0_2_2_out ),
       .io_V_wire_in_33( VwireModule_io_VwirePorts_0_2_1_out ),
       .io_V_wire_in_32( VwireModule_io_VwirePorts_0_2_0_out ),
       .io_V_wire_in_31( VwireModule_io_VwirePorts_0_1_15_out ),
       .io_V_wire_in_30( VwireModule_io_VwirePorts_0_1_14_out ),
       .io_V_wire_in_29( VwireModule_io_VwirePorts_0_1_13_out ),
       .io_V_wire_in_28( VwireModule_io_VwirePorts_0_1_12_out ),
       .io_V_wire_in_27( VwireModule_io_VwirePorts_0_1_11_out ),
       .io_V_wire_in_26( VwireModule_io_VwirePorts_0_1_10_out ),
       .io_V_wire_in_25( VwireModule_io_VwirePorts_0_1_9_out ),
       .io_V_wire_in_24( VwireModule_io_VwirePorts_0_1_8_out ),
       .io_V_wire_in_23( VwireModule_io_VwirePorts_0_1_7_out ),
       .io_V_wire_in_22( VwireModule_io_VwirePorts_0_1_6_out ),
       .io_V_wire_in_21( VwireModule_io_VwirePorts_0_1_5_out ),
       .io_V_wire_in_20( VwireModule_io_VwirePorts_0_1_4_out ),
       .io_V_wire_in_19( VwireModule_io_VwirePorts_0_1_3_out ),
       .io_V_wire_in_18( VwireModule_io_VwirePorts_0_1_2_out ),
       .io_V_wire_in_17( VwireModule_io_VwirePorts_0_1_1_out ),
       .io_V_wire_in_16( VwireModule_io_VwirePorts_0_1_0_out ),
       .io_V_wire_in_15( VwireModule_io_VwirePorts_0_0_15_out ),
       .io_V_wire_in_14( VwireModule_io_VwirePorts_0_0_14_out ),
       .io_V_wire_in_13( VwireModule_io_VwirePorts_0_0_13_out ),
       .io_V_wire_in_12( VwireModule_io_VwirePorts_0_0_12_out ),
       .io_V_wire_in_11( VwireModule_io_VwirePorts_0_0_11_out ),
       .io_V_wire_in_10( VwireModule_io_VwirePorts_0_0_10_out ),
       .io_V_wire_in_9( VwireModule_io_VwirePorts_0_0_9_out ),
       .io_V_wire_in_8( VwireModule_io_VwirePorts_0_0_8_out ),
       .io_V_wire_in_7( VwireModule_io_VwirePorts_0_0_7_out ),
       .io_V_wire_in_6( VwireModule_io_VwirePorts_0_0_6_out ),
       .io_V_wire_in_5( VwireModule_io_VwirePorts_0_0_5_out ),
       .io_V_wire_in_4( VwireModule_io_VwirePorts_0_0_4_out ),
       .io_V_wire_in_3( VwireModule_io_VwirePorts_0_0_3_out ),
       .io_V_wire_in_2( VwireModule_io_VwirePorts_0_0_2_out ),
       .io_V_wire_in_1( VwireModule_io_VwirePorts_0_0_1_out ),
       .io_V_wire_in_0( VwireModule_io_VwirePorts_0_0_0_out ),
       .io_V_wire_out_367( ArrayRowModule_io_V_wire_out_367 ),
       .io_V_wire_out_366( ArrayRowModule_io_V_wire_out_366 ),
       .io_V_wire_out_365( ArrayRowModule_io_V_wire_out_365 ),
       .io_V_wire_out_364( ArrayRowModule_io_V_wire_out_364 ),
       .io_V_wire_out_363( ArrayRowModule_io_V_wire_out_363 ),
       .io_V_wire_out_362( ArrayRowModule_io_V_wire_out_362 ),
       .io_V_wire_out_361( ArrayRowModule_io_V_wire_out_361 ),
       .io_V_wire_out_360( ArrayRowModule_io_V_wire_out_360 ),
       .io_V_wire_out_359( ArrayRowModule_io_V_wire_out_359 ),
       .io_V_wire_out_358( ArrayRowModule_io_V_wire_out_358 ),
       .io_V_wire_out_357( ArrayRowModule_io_V_wire_out_357 ),
       .io_V_wire_out_356( ArrayRowModule_io_V_wire_out_356 ),
       .io_V_wire_out_355( ArrayRowModule_io_V_wire_out_355 ),
       .io_V_wire_out_354( ArrayRowModule_io_V_wire_out_354 ),
       .io_V_wire_out_353( ArrayRowModule_io_V_wire_out_353 ),
       .io_V_wire_out_352( ArrayRowModule_io_V_wire_out_352 ),
       .io_V_wire_out_351( ArrayRowModule_io_V_wire_out_351 ),
       .io_V_wire_out_350( ArrayRowModule_io_V_wire_out_350 ),
       .io_V_wire_out_349( ArrayRowModule_io_V_wire_out_349 ),
       .io_V_wire_out_348( ArrayRowModule_io_V_wire_out_348 ),
       .io_V_wire_out_347( ArrayRowModule_io_V_wire_out_347 ),
       .io_V_wire_out_346( ArrayRowModule_io_V_wire_out_346 ),
       .io_V_wire_out_345( ArrayRowModule_io_V_wire_out_345 ),
       .io_V_wire_out_344( ArrayRowModule_io_V_wire_out_344 ),
       .io_V_wire_out_343( ArrayRowModule_io_V_wire_out_343 ),
       .io_V_wire_out_342( ArrayRowModule_io_V_wire_out_342 ),
       .io_V_wire_out_341( ArrayRowModule_io_V_wire_out_341 ),
       .io_V_wire_out_340( ArrayRowModule_io_V_wire_out_340 ),
       .io_V_wire_out_339( ArrayRowModule_io_V_wire_out_339 ),
       .io_V_wire_out_338( ArrayRowModule_io_V_wire_out_338 ),
       .io_V_wire_out_337( ArrayRowModule_io_V_wire_out_337 ),
       .io_V_wire_out_336( ArrayRowModule_io_V_wire_out_336 ),
       .io_V_wire_out_335( ArrayRowModule_io_V_wire_out_335 ),
       .io_V_wire_out_334( ArrayRowModule_io_V_wire_out_334 ),
       .io_V_wire_out_333( ArrayRowModule_io_V_wire_out_333 ),
       .io_V_wire_out_332( ArrayRowModule_io_V_wire_out_332 ),
       .io_V_wire_out_331( ArrayRowModule_io_V_wire_out_331 ),
       .io_V_wire_out_330( ArrayRowModule_io_V_wire_out_330 ),
       .io_V_wire_out_329( ArrayRowModule_io_V_wire_out_329 ),
       .io_V_wire_out_328( ArrayRowModule_io_V_wire_out_328 ),
       .io_V_wire_out_327( ArrayRowModule_io_V_wire_out_327 ),
       .io_V_wire_out_326( ArrayRowModule_io_V_wire_out_326 ),
       .io_V_wire_out_325( ArrayRowModule_io_V_wire_out_325 ),
       .io_V_wire_out_324( ArrayRowModule_io_V_wire_out_324 ),
       .io_V_wire_out_323( ArrayRowModule_io_V_wire_out_323 ),
       .io_V_wire_out_322( ArrayRowModule_io_V_wire_out_322 ),
       .io_V_wire_out_321( ArrayRowModule_io_V_wire_out_321 ),
       .io_V_wire_out_320( ArrayRowModule_io_V_wire_out_320 ),
       .io_V_wire_out_319( ArrayRowModule_io_V_wire_out_319 ),
       .io_V_wire_out_318( ArrayRowModule_io_V_wire_out_318 ),
       .io_V_wire_out_317( ArrayRowModule_io_V_wire_out_317 ),
       .io_V_wire_out_316( ArrayRowModule_io_V_wire_out_316 ),
       .io_V_wire_out_315( ArrayRowModule_io_V_wire_out_315 ),
       .io_V_wire_out_314( ArrayRowModule_io_V_wire_out_314 ),
       .io_V_wire_out_313( ArrayRowModule_io_V_wire_out_313 ),
       .io_V_wire_out_312( ArrayRowModule_io_V_wire_out_312 ),
       .io_V_wire_out_311( ArrayRowModule_io_V_wire_out_311 ),
       .io_V_wire_out_310( ArrayRowModule_io_V_wire_out_310 ),
       .io_V_wire_out_309( ArrayRowModule_io_V_wire_out_309 ),
       .io_V_wire_out_308( ArrayRowModule_io_V_wire_out_308 ),
       .io_V_wire_out_307( ArrayRowModule_io_V_wire_out_307 ),
       .io_V_wire_out_306( ArrayRowModule_io_V_wire_out_306 ),
       .io_V_wire_out_305( ArrayRowModule_io_V_wire_out_305 ),
       .io_V_wire_out_304( ArrayRowModule_io_V_wire_out_304 ),
       .io_V_wire_out_303( ArrayRowModule_io_V_wire_out_303 ),
       .io_V_wire_out_302( ArrayRowModule_io_V_wire_out_302 ),
       .io_V_wire_out_301( ArrayRowModule_io_V_wire_out_301 ),
       .io_V_wire_out_300( ArrayRowModule_io_V_wire_out_300 ),
       .io_V_wire_out_299( ArrayRowModule_io_V_wire_out_299 ),
       .io_V_wire_out_298( ArrayRowModule_io_V_wire_out_298 ),
       .io_V_wire_out_297( ArrayRowModule_io_V_wire_out_297 ),
       .io_V_wire_out_296( ArrayRowModule_io_V_wire_out_296 ),
       .io_V_wire_out_295( ArrayRowModule_io_V_wire_out_295 ),
       .io_V_wire_out_294( ArrayRowModule_io_V_wire_out_294 ),
       .io_V_wire_out_293( ArrayRowModule_io_V_wire_out_293 ),
       .io_V_wire_out_292( ArrayRowModule_io_V_wire_out_292 ),
       .io_V_wire_out_291( ArrayRowModule_io_V_wire_out_291 ),
       .io_V_wire_out_290( ArrayRowModule_io_V_wire_out_290 ),
       .io_V_wire_out_289( ArrayRowModule_io_V_wire_out_289 ),
       .io_V_wire_out_288( ArrayRowModule_io_V_wire_out_288 ),
       .io_V_wire_out_287( ArrayRowModule_io_V_wire_out_287 ),
       .io_V_wire_out_286( ArrayRowModule_io_V_wire_out_286 ),
       .io_V_wire_out_285( ArrayRowModule_io_V_wire_out_285 ),
       .io_V_wire_out_284( ArrayRowModule_io_V_wire_out_284 ),
       .io_V_wire_out_283( ArrayRowModule_io_V_wire_out_283 ),
       .io_V_wire_out_282( ArrayRowModule_io_V_wire_out_282 ),
       .io_V_wire_out_281( ArrayRowModule_io_V_wire_out_281 ),
       .io_V_wire_out_280( ArrayRowModule_io_V_wire_out_280 ),
       .io_V_wire_out_279( ArrayRowModule_io_V_wire_out_279 ),
       .io_V_wire_out_278( ArrayRowModule_io_V_wire_out_278 ),
       .io_V_wire_out_277( ArrayRowModule_io_V_wire_out_277 ),
       .io_V_wire_out_276( ArrayRowModule_io_V_wire_out_276 ),
       .io_V_wire_out_275( ArrayRowModule_io_V_wire_out_275 ),
       .io_V_wire_out_274( ArrayRowModule_io_V_wire_out_274 ),
       .io_V_wire_out_273( ArrayRowModule_io_V_wire_out_273 ),
       .io_V_wire_out_272( ArrayRowModule_io_V_wire_out_272 ),
       .io_V_wire_out_271( ArrayRowModule_io_V_wire_out_271 ),
       .io_V_wire_out_270( ArrayRowModule_io_V_wire_out_270 ),
       .io_V_wire_out_269( ArrayRowModule_io_V_wire_out_269 ),
       .io_V_wire_out_268( ArrayRowModule_io_V_wire_out_268 ),
       .io_V_wire_out_267( ArrayRowModule_io_V_wire_out_267 ),
       .io_V_wire_out_266( ArrayRowModule_io_V_wire_out_266 ),
       .io_V_wire_out_265( ArrayRowModule_io_V_wire_out_265 ),
       .io_V_wire_out_264( ArrayRowModule_io_V_wire_out_264 ),
       .io_V_wire_out_263( ArrayRowModule_io_V_wire_out_263 ),
       .io_V_wire_out_262( ArrayRowModule_io_V_wire_out_262 ),
       .io_V_wire_out_261( ArrayRowModule_io_V_wire_out_261 ),
       .io_V_wire_out_260( ArrayRowModule_io_V_wire_out_260 ),
       .io_V_wire_out_259( ArrayRowModule_io_V_wire_out_259 ),
       .io_V_wire_out_258( ArrayRowModule_io_V_wire_out_258 ),
       .io_V_wire_out_257( ArrayRowModule_io_V_wire_out_257 ),
       .io_V_wire_out_256( ArrayRowModule_io_V_wire_out_256 ),
       .io_V_wire_out_255( ArrayRowModule_io_V_wire_out_255 ),
       .io_V_wire_out_254( ArrayRowModule_io_V_wire_out_254 ),
       .io_V_wire_out_253( ArrayRowModule_io_V_wire_out_253 ),
       .io_V_wire_out_252( ArrayRowModule_io_V_wire_out_252 ),
       .io_V_wire_out_251( ArrayRowModule_io_V_wire_out_251 ),
       .io_V_wire_out_250( ArrayRowModule_io_V_wire_out_250 ),
       .io_V_wire_out_249( ArrayRowModule_io_V_wire_out_249 ),
       .io_V_wire_out_248( ArrayRowModule_io_V_wire_out_248 ),
       .io_V_wire_out_247( ArrayRowModule_io_V_wire_out_247 ),
       .io_V_wire_out_246( ArrayRowModule_io_V_wire_out_246 ),
       .io_V_wire_out_245( ArrayRowModule_io_V_wire_out_245 ),
       .io_V_wire_out_244( ArrayRowModule_io_V_wire_out_244 ),
       .io_V_wire_out_243( ArrayRowModule_io_V_wire_out_243 ),
       .io_V_wire_out_242( ArrayRowModule_io_V_wire_out_242 ),
       .io_V_wire_out_241( ArrayRowModule_io_V_wire_out_241 ),
       .io_V_wire_out_240( ArrayRowModule_io_V_wire_out_240 ),
       .io_V_wire_out_239( ArrayRowModule_io_V_wire_out_239 ),
       .io_V_wire_out_238( ArrayRowModule_io_V_wire_out_238 ),
       .io_V_wire_out_237( ArrayRowModule_io_V_wire_out_237 ),
       .io_V_wire_out_236( ArrayRowModule_io_V_wire_out_236 ),
       .io_V_wire_out_235( ArrayRowModule_io_V_wire_out_235 ),
       .io_V_wire_out_234( ArrayRowModule_io_V_wire_out_234 ),
       .io_V_wire_out_233( ArrayRowModule_io_V_wire_out_233 ),
       .io_V_wire_out_232( ArrayRowModule_io_V_wire_out_232 ),
       .io_V_wire_out_231( ArrayRowModule_io_V_wire_out_231 ),
       .io_V_wire_out_230( ArrayRowModule_io_V_wire_out_230 ),
       .io_V_wire_out_229( ArrayRowModule_io_V_wire_out_229 ),
       .io_V_wire_out_228( ArrayRowModule_io_V_wire_out_228 ),
       .io_V_wire_out_227( ArrayRowModule_io_V_wire_out_227 ),
       .io_V_wire_out_226( ArrayRowModule_io_V_wire_out_226 ),
       .io_V_wire_out_225( ArrayRowModule_io_V_wire_out_225 ),
       .io_V_wire_out_224( ArrayRowModule_io_V_wire_out_224 ),
       .io_V_wire_out_223( ArrayRowModule_io_V_wire_out_223 ),
       .io_V_wire_out_222( ArrayRowModule_io_V_wire_out_222 ),
       .io_V_wire_out_221( ArrayRowModule_io_V_wire_out_221 ),
       .io_V_wire_out_220( ArrayRowModule_io_V_wire_out_220 ),
       .io_V_wire_out_219( ArrayRowModule_io_V_wire_out_219 ),
       .io_V_wire_out_218( ArrayRowModule_io_V_wire_out_218 ),
       .io_V_wire_out_217( ArrayRowModule_io_V_wire_out_217 ),
       .io_V_wire_out_216( ArrayRowModule_io_V_wire_out_216 ),
       .io_V_wire_out_215( ArrayRowModule_io_V_wire_out_215 ),
       .io_V_wire_out_214( ArrayRowModule_io_V_wire_out_214 ),
       .io_V_wire_out_213( ArrayRowModule_io_V_wire_out_213 ),
       .io_V_wire_out_212( ArrayRowModule_io_V_wire_out_212 ),
       .io_V_wire_out_211( ArrayRowModule_io_V_wire_out_211 ),
       .io_V_wire_out_210( ArrayRowModule_io_V_wire_out_210 ),
       .io_V_wire_out_209( ArrayRowModule_io_V_wire_out_209 ),
       .io_V_wire_out_208( ArrayRowModule_io_V_wire_out_208 ),
       .io_V_wire_out_207( ArrayRowModule_io_V_wire_out_207 ),
       .io_V_wire_out_206( ArrayRowModule_io_V_wire_out_206 ),
       .io_V_wire_out_205( ArrayRowModule_io_V_wire_out_205 ),
       .io_V_wire_out_204( ArrayRowModule_io_V_wire_out_204 ),
       .io_V_wire_out_203( ArrayRowModule_io_V_wire_out_203 ),
       .io_V_wire_out_202( ArrayRowModule_io_V_wire_out_202 ),
       .io_V_wire_out_201( ArrayRowModule_io_V_wire_out_201 ),
       .io_V_wire_out_200( ArrayRowModule_io_V_wire_out_200 ),
       .io_V_wire_out_199( ArrayRowModule_io_V_wire_out_199 ),
       .io_V_wire_out_198( ArrayRowModule_io_V_wire_out_198 ),
       .io_V_wire_out_197( ArrayRowModule_io_V_wire_out_197 ),
       .io_V_wire_out_196( ArrayRowModule_io_V_wire_out_196 ),
       .io_V_wire_out_195( ArrayRowModule_io_V_wire_out_195 ),
       .io_V_wire_out_194( ArrayRowModule_io_V_wire_out_194 ),
       .io_V_wire_out_193( ArrayRowModule_io_V_wire_out_193 ),
       .io_V_wire_out_192( ArrayRowModule_io_V_wire_out_192 ),
       .io_V_wire_out_191( ArrayRowModule_io_V_wire_out_191 ),
       .io_V_wire_out_190( ArrayRowModule_io_V_wire_out_190 ),
       .io_V_wire_out_189( ArrayRowModule_io_V_wire_out_189 ),
       .io_V_wire_out_188( ArrayRowModule_io_V_wire_out_188 ),
       .io_V_wire_out_187( ArrayRowModule_io_V_wire_out_187 ),
       .io_V_wire_out_186( ArrayRowModule_io_V_wire_out_186 ),
       .io_V_wire_out_185( ArrayRowModule_io_V_wire_out_185 ),
       .io_V_wire_out_184( ArrayRowModule_io_V_wire_out_184 ),
       .io_V_wire_out_183( ArrayRowModule_io_V_wire_out_183 ),
       .io_V_wire_out_182( ArrayRowModule_io_V_wire_out_182 ),
       .io_V_wire_out_181( ArrayRowModule_io_V_wire_out_181 ),
       .io_V_wire_out_180( ArrayRowModule_io_V_wire_out_180 ),
       .io_V_wire_out_179( ArrayRowModule_io_V_wire_out_179 ),
       .io_V_wire_out_178( ArrayRowModule_io_V_wire_out_178 ),
       .io_V_wire_out_177( ArrayRowModule_io_V_wire_out_177 ),
       .io_V_wire_out_176( ArrayRowModule_io_V_wire_out_176 ),
       .io_V_wire_out_175( ArrayRowModule_io_V_wire_out_175 ),
       .io_V_wire_out_174( ArrayRowModule_io_V_wire_out_174 ),
       .io_V_wire_out_173( ArrayRowModule_io_V_wire_out_173 ),
       .io_V_wire_out_172( ArrayRowModule_io_V_wire_out_172 ),
       .io_V_wire_out_171( ArrayRowModule_io_V_wire_out_171 ),
       .io_V_wire_out_170( ArrayRowModule_io_V_wire_out_170 ),
       .io_V_wire_out_169( ArrayRowModule_io_V_wire_out_169 ),
       .io_V_wire_out_168( ArrayRowModule_io_V_wire_out_168 ),
       .io_V_wire_out_167( ArrayRowModule_io_V_wire_out_167 ),
       .io_V_wire_out_166( ArrayRowModule_io_V_wire_out_166 ),
       .io_V_wire_out_165( ArrayRowModule_io_V_wire_out_165 ),
       .io_V_wire_out_164( ArrayRowModule_io_V_wire_out_164 ),
       .io_V_wire_out_163( ArrayRowModule_io_V_wire_out_163 ),
       .io_V_wire_out_162( ArrayRowModule_io_V_wire_out_162 ),
       .io_V_wire_out_161( ArrayRowModule_io_V_wire_out_161 ),
       .io_V_wire_out_160( ArrayRowModule_io_V_wire_out_160 ),
       .io_V_wire_out_159( ArrayRowModule_io_V_wire_out_159 ),
       .io_V_wire_out_158( ArrayRowModule_io_V_wire_out_158 ),
       .io_V_wire_out_157( ArrayRowModule_io_V_wire_out_157 ),
       .io_V_wire_out_156( ArrayRowModule_io_V_wire_out_156 ),
       .io_V_wire_out_155( ArrayRowModule_io_V_wire_out_155 ),
       .io_V_wire_out_154( ArrayRowModule_io_V_wire_out_154 ),
       .io_V_wire_out_153( ArrayRowModule_io_V_wire_out_153 ),
       .io_V_wire_out_152( ArrayRowModule_io_V_wire_out_152 ),
       .io_V_wire_out_151( ArrayRowModule_io_V_wire_out_151 ),
       .io_V_wire_out_150( ArrayRowModule_io_V_wire_out_150 ),
       .io_V_wire_out_149( ArrayRowModule_io_V_wire_out_149 ),
       .io_V_wire_out_148( ArrayRowModule_io_V_wire_out_148 ),
       .io_V_wire_out_147( ArrayRowModule_io_V_wire_out_147 ),
       .io_V_wire_out_146( ArrayRowModule_io_V_wire_out_146 ),
       .io_V_wire_out_145( ArrayRowModule_io_V_wire_out_145 ),
       .io_V_wire_out_144( ArrayRowModule_io_V_wire_out_144 ),
       .io_V_wire_out_143( ArrayRowModule_io_V_wire_out_143 ),
       .io_V_wire_out_142( ArrayRowModule_io_V_wire_out_142 ),
       .io_V_wire_out_141( ArrayRowModule_io_V_wire_out_141 ),
       .io_V_wire_out_140( ArrayRowModule_io_V_wire_out_140 ),
       .io_V_wire_out_139( ArrayRowModule_io_V_wire_out_139 ),
       .io_V_wire_out_138( ArrayRowModule_io_V_wire_out_138 ),
       .io_V_wire_out_137( ArrayRowModule_io_V_wire_out_137 ),
       .io_V_wire_out_136( ArrayRowModule_io_V_wire_out_136 ),
       .io_V_wire_out_135( ArrayRowModule_io_V_wire_out_135 ),
       .io_V_wire_out_134( ArrayRowModule_io_V_wire_out_134 ),
       .io_V_wire_out_133( ArrayRowModule_io_V_wire_out_133 ),
       .io_V_wire_out_132( ArrayRowModule_io_V_wire_out_132 ),
       .io_V_wire_out_131( ArrayRowModule_io_V_wire_out_131 ),
       .io_V_wire_out_130( ArrayRowModule_io_V_wire_out_130 ),
       .io_V_wire_out_129( ArrayRowModule_io_V_wire_out_129 ),
       .io_V_wire_out_128( ArrayRowModule_io_V_wire_out_128 ),
       .io_V_wire_out_127( ArrayRowModule_io_V_wire_out_127 ),
       .io_V_wire_out_126( ArrayRowModule_io_V_wire_out_126 ),
       .io_V_wire_out_125( ArrayRowModule_io_V_wire_out_125 ),
       .io_V_wire_out_124( ArrayRowModule_io_V_wire_out_124 ),
       .io_V_wire_out_123( ArrayRowModule_io_V_wire_out_123 ),
       .io_V_wire_out_122( ArrayRowModule_io_V_wire_out_122 ),
       .io_V_wire_out_121( ArrayRowModule_io_V_wire_out_121 ),
       .io_V_wire_out_120( ArrayRowModule_io_V_wire_out_120 ),
       .io_V_wire_out_119( ArrayRowModule_io_V_wire_out_119 ),
       .io_V_wire_out_118( ArrayRowModule_io_V_wire_out_118 ),
       .io_V_wire_out_117( ArrayRowModule_io_V_wire_out_117 ),
       .io_V_wire_out_116( ArrayRowModule_io_V_wire_out_116 ),
       .io_V_wire_out_115( ArrayRowModule_io_V_wire_out_115 ),
       .io_V_wire_out_114( ArrayRowModule_io_V_wire_out_114 ),
       .io_V_wire_out_113( ArrayRowModule_io_V_wire_out_113 ),
       .io_V_wire_out_112( ArrayRowModule_io_V_wire_out_112 ),
       .io_V_wire_out_111( ArrayRowModule_io_V_wire_out_111 ),
       .io_V_wire_out_110( ArrayRowModule_io_V_wire_out_110 ),
       .io_V_wire_out_109( ArrayRowModule_io_V_wire_out_109 ),
       .io_V_wire_out_108( ArrayRowModule_io_V_wire_out_108 ),
       .io_V_wire_out_107( ArrayRowModule_io_V_wire_out_107 ),
       .io_V_wire_out_106( ArrayRowModule_io_V_wire_out_106 ),
       .io_V_wire_out_105( ArrayRowModule_io_V_wire_out_105 ),
       .io_V_wire_out_104( ArrayRowModule_io_V_wire_out_104 ),
       .io_V_wire_out_103( ArrayRowModule_io_V_wire_out_103 ),
       .io_V_wire_out_102( ArrayRowModule_io_V_wire_out_102 ),
       .io_V_wire_out_101( ArrayRowModule_io_V_wire_out_101 ),
       .io_V_wire_out_100( ArrayRowModule_io_V_wire_out_100 ),
       .io_V_wire_out_99( ArrayRowModule_io_V_wire_out_99 ),
       .io_V_wire_out_98( ArrayRowModule_io_V_wire_out_98 ),
       .io_V_wire_out_97( ArrayRowModule_io_V_wire_out_97 ),
       .io_V_wire_out_96( ArrayRowModule_io_V_wire_out_96 ),
       .io_V_wire_out_95( ArrayRowModule_io_V_wire_out_95 ),
       .io_V_wire_out_94( ArrayRowModule_io_V_wire_out_94 ),
       .io_V_wire_out_93( ArrayRowModule_io_V_wire_out_93 ),
       .io_V_wire_out_92( ArrayRowModule_io_V_wire_out_92 ),
       .io_V_wire_out_91( ArrayRowModule_io_V_wire_out_91 ),
       .io_V_wire_out_90( ArrayRowModule_io_V_wire_out_90 ),
       .io_V_wire_out_89( ArrayRowModule_io_V_wire_out_89 ),
       .io_V_wire_out_88( ArrayRowModule_io_V_wire_out_88 ),
       .io_V_wire_out_87( ArrayRowModule_io_V_wire_out_87 ),
       .io_V_wire_out_86( ArrayRowModule_io_V_wire_out_86 ),
       .io_V_wire_out_85( ArrayRowModule_io_V_wire_out_85 ),
       .io_V_wire_out_84( ArrayRowModule_io_V_wire_out_84 ),
       .io_V_wire_out_83( ArrayRowModule_io_V_wire_out_83 ),
       .io_V_wire_out_82( ArrayRowModule_io_V_wire_out_82 ),
       .io_V_wire_out_81( ArrayRowModule_io_V_wire_out_81 ),
       .io_V_wire_out_80( ArrayRowModule_io_V_wire_out_80 ),
       .io_V_wire_out_79( ArrayRowModule_io_V_wire_out_79 ),
       .io_V_wire_out_78( ArrayRowModule_io_V_wire_out_78 ),
       .io_V_wire_out_77( ArrayRowModule_io_V_wire_out_77 ),
       .io_V_wire_out_76( ArrayRowModule_io_V_wire_out_76 ),
       .io_V_wire_out_75( ArrayRowModule_io_V_wire_out_75 ),
       .io_V_wire_out_74( ArrayRowModule_io_V_wire_out_74 ),
       .io_V_wire_out_73( ArrayRowModule_io_V_wire_out_73 ),
       .io_V_wire_out_72( ArrayRowModule_io_V_wire_out_72 ),
       .io_V_wire_out_71( ArrayRowModule_io_V_wire_out_71 ),
       .io_V_wire_out_70( ArrayRowModule_io_V_wire_out_70 ),
       .io_V_wire_out_69( ArrayRowModule_io_V_wire_out_69 ),
       .io_V_wire_out_68( ArrayRowModule_io_V_wire_out_68 ),
       .io_V_wire_out_67( ArrayRowModule_io_V_wire_out_67 ),
       .io_V_wire_out_66( ArrayRowModule_io_V_wire_out_66 ),
       .io_V_wire_out_65( ArrayRowModule_io_V_wire_out_65 ),
       .io_V_wire_out_64( ArrayRowModule_io_V_wire_out_64 ),
       .io_V_wire_out_63( ArrayRowModule_io_V_wire_out_63 ),
       .io_V_wire_out_62( ArrayRowModule_io_V_wire_out_62 ),
       .io_V_wire_out_61( ArrayRowModule_io_V_wire_out_61 ),
       .io_V_wire_out_60( ArrayRowModule_io_V_wire_out_60 ),
       .io_V_wire_out_59( ArrayRowModule_io_V_wire_out_59 ),
       .io_V_wire_out_58( ArrayRowModule_io_V_wire_out_58 ),
       .io_V_wire_out_57( ArrayRowModule_io_V_wire_out_57 ),
       .io_V_wire_out_56( ArrayRowModule_io_V_wire_out_56 ),
       .io_V_wire_out_55( ArrayRowModule_io_V_wire_out_55 ),
       .io_V_wire_out_54( ArrayRowModule_io_V_wire_out_54 ),
       .io_V_wire_out_53( ArrayRowModule_io_V_wire_out_53 ),
       .io_V_wire_out_52( ArrayRowModule_io_V_wire_out_52 ),
       .io_V_wire_out_51( ArrayRowModule_io_V_wire_out_51 ),
       .io_V_wire_out_50( ArrayRowModule_io_V_wire_out_50 ),
       .io_V_wire_out_49( ArrayRowModule_io_V_wire_out_49 ),
       .io_V_wire_out_48( ArrayRowModule_io_V_wire_out_48 ),
       .io_V_wire_out_47( ArrayRowModule_io_V_wire_out_47 ),
       .io_V_wire_out_46( ArrayRowModule_io_V_wire_out_46 ),
       .io_V_wire_out_45( ArrayRowModule_io_V_wire_out_45 ),
       .io_V_wire_out_44( ArrayRowModule_io_V_wire_out_44 ),
       .io_V_wire_out_43( ArrayRowModule_io_V_wire_out_43 ),
       .io_V_wire_out_42( ArrayRowModule_io_V_wire_out_42 ),
       .io_V_wire_out_41( ArrayRowModule_io_V_wire_out_41 ),
       .io_V_wire_out_40( ArrayRowModule_io_V_wire_out_40 ),
       .io_V_wire_out_39( ArrayRowModule_io_V_wire_out_39 ),
       .io_V_wire_out_38( ArrayRowModule_io_V_wire_out_38 ),
       .io_V_wire_out_37( ArrayRowModule_io_V_wire_out_37 ),
       .io_V_wire_out_36( ArrayRowModule_io_V_wire_out_36 ),
       .io_V_wire_out_35( ArrayRowModule_io_V_wire_out_35 ),
       .io_V_wire_out_34( ArrayRowModule_io_V_wire_out_34 ),
       .io_V_wire_out_33( ArrayRowModule_io_V_wire_out_33 ),
       .io_V_wire_out_32( ArrayRowModule_io_V_wire_out_32 ),
       .io_V_wire_out_31( ArrayRowModule_io_V_wire_out_31 ),
       .io_V_wire_out_30( ArrayRowModule_io_V_wire_out_30 ),
       .io_V_wire_out_29( ArrayRowModule_io_V_wire_out_29 ),
       .io_V_wire_out_28( ArrayRowModule_io_V_wire_out_28 ),
       .io_V_wire_out_27( ArrayRowModule_io_V_wire_out_27 ),
       .io_V_wire_out_26( ArrayRowModule_io_V_wire_out_26 ),
       .io_V_wire_out_25( ArrayRowModule_io_V_wire_out_25 ),
       .io_V_wire_out_24( ArrayRowModule_io_V_wire_out_24 ),
       .io_V_wire_out_23( ArrayRowModule_io_V_wire_out_23 ),
       .io_V_wire_out_22( ArrayRowModule_io_V_wire_out_22 ),
       .io_V_wire_out_21( ArrayRowModule_io_V_wire_out_21 ),
       .io_V_wire_out_20( ArrayRowModule_io_V_wire_out_20 ),
       .io_V_wire_out_19( ArrayRowModule_io_V_wire_out_19 ),
       .io_V_wire_out_18( ArrayRowModule_io_V_wire_out_18 ),
       .io_V_wire_out_17( ArrayRowModule_io_V_wire_out_17 ),
       .io_V_wire_out_16( ArrayRowModule_io_V_wire_out_16 ),
       .io_V_wire_out_15( ArrayRowModule_io_V_wire_out_15 ),
       .io_V_wire_out_14( ArrayRowModule_io_V_wire_out_14 ),
       .io_V_wire_out_13( ArrayRowModule_io_V_wire_out_13 ),
       .io_V_wire_out_12( ArrayRowModule_io_V_wire_out_12 ),
       .io_V_wire_out_11( ArrayRowModule_io_V_wire_out_11 ),
       .io_V_wire_out_10( ArrayRowModule_io_V_wire_out_10 ),
       .io_V_wire_out_9( ArrayRowModule_io_V_wire_out_9 ),
       .io_V_wire_out_8( ArrayRowModule_io_V_wire_out_8 ),
       .io_V_wire_out_7( ArrayRowModule_io_V_wire_out_7 ),
       .io_V_wire_out_6( ArrayRowModule_io_V_wire_out_6 ),
       .io_V_wire_out_5( ArrayRowModule_io_V_wire_out_5 ),
       .io_V_wire_out_4( ArrayRowModule_io_V_wire_out_4 ),
       .io_V_wire_out_3( ArrayRowModule_io_V_wire_out_3 ),
       .io_V_wire_out_2( ArrayRowModule_io_V_wire_out_2 ),
       .io_V_wire_out_1( ArrayRowModule_io_V_wire_out_1 ),
       .io_V_wire_out_0( ArrayRowModule_io_V_wire_out_0 ),
       .io_V_wire_en_22( ArrayRowModule_io_V_wire_en_22 ),
       .io_V_wire_en_21( ArrayRowModule_io_V_wire_en_21 ),
       .io_V_wire_en_20( ArrayRowModule_io_V_wire_en_20 ),
       .io_V_wire_en_19( ArrayRowModule_io_V_wire_en_19 ),
       .io_V_wire_en_18( ArrayRowModule_io_V_wire_en_18 ),
       .io_V_wire_en_17( ArrayRowModule_io_V_wire_en_17 ),
       .io_V_wire_en_16( ArrayRowModule_io_V_wire_en_16 ),
       .io_V_wire_en_15( ArrayRowModule_io_V_wire_en_15 ),
       .io_V_wire_en_14( ArrayRowModule_io_V_wire_en_14 ),
       .io_V_wire_en_13( ArrayRowModule_io_V_wire_en_13 ),
       .io_V_wire_en_12( ArrayRowModule_io_V_wire_en_12 ),
       .io_V_wire_en_11( ArrayRowModule_io_V_wire_en_11 ),
       .io_V_wire_en_10( ArrayRowModule_io_V_wire_en_10 ),
       .io_V_wire_en_9( ArrayRowModule_io_V_wire_en_9 ),
       .io_V_wire_en_8( ArrayRowModule_io_V_wire_en_8 ),
       .io_V_wire_en_7( ArrayRowModule_io_V_wire_en_7 ),
       .io_V_wire_en_6( ArrayRowModule_io_V_wire_en_6 ),
       .io_V_wire_en_5( ArrayRowModule_io_V_wire_en_5 ),
       .io_V_wire_en_4( ArrayRowModule_io_V_wire_en_4 ),
       .io_V_wire_en_3( ArrayRowModule_io_V_wire_en_3 ),
       .io_V_wire_en_2( ArrayRowModule_io_V_wire_en_2 ),
       .io_V_wire_en_1( ArrayRowModule_io_V_wire_en_1 ),
       .io_V_wire_en_0( ArrayRowModule_io_V_wire_en_0 ),
       .io_G_wire_above_3( T1535 ),
       .io_G_wire_above_2( T1534 ),
       .io_G_wire_above_1( T1533 ),
       .io_G_wire_above_0( T1532 ),
       .io_H_wire_above_32( T1531 ),
       .io_H_wire_above_31( T1530 ),
       .io_H_wire_above_30( T1529 ),
       .io_H_wire_above_29( T1528 ),
       .io_H_wire_above_28( T1527 ),
       .io_H_wire_above_27( T1526 ),
       .io_H_wire_above_26( T1525 ),
       .io_H_wire_above_25( T1524 ),
       .io_H_wire_above_24( T1523 ),
       .io_H_wire_above_23( T1522 ),
       .io_H_wire_above_22( T1521 ),
       .io_H_wire_above_21( T1520 ),
       .io_H_wire_above_20( T1519 ),
       .io_H_wire_above_19( T1518 ),
       .io_H_wire_above_18( T1517 ),
       .io_H_wire_above_17( T1516 ),
       .io_H_wire_above_16( T1515 ),
       .io_H_wire_above_15( T1514 ),
       .io_H_wire_above_14( T1513 ),
       .io_H_wire_above_13( T1512 ),
       .io_H_wire_above_12( T1511 ),
       .io_H_wire_above_11( T1510 ),
       .io_H_wire_above_10( T1509 ),
       .io_H_wire_above_9( T1508 ),
       .io_H_wire_above_8( T1507 ),
       .io_H_wire_above_7( T1506 ),
       .io_H_wire_above_6( T1505 ),
       .io_H_wire_above_5( T1504 ),
       .io_H_wire_above_4( T1503 ),
       .io_H_wire_above_3( T1502 ),
       .io_H_wire_above_2( T1501 ),
       .io_H_wire_above_1( T1500 ),
       .io_H_wire_above_0( T1499 ),
       .io_mem_bus_in_23( io_mem_bus_in_23 ),
       .io_mem_bus_in_22( io_mem_bus_in_22 ),
       .io_mem_bus_in_21( io_mem_bus_in_21 ),
       .io_mem_bus_in_20( io_mem_bus_in_20 ),
       .io_mem_bus_in_19( io_mem_bus_in_19 ),
       .io_mem_bus_in_18( io_mem_bus_in_18 ),
       .io_mem_bus_in_17( io_mem_bus_in_17 ),
       .io_mem_bus_in_16( io_mem_bus_in_16 ),
       .io_mem_bus_in_15( io_mem_bus_in_15 ),
       .io_mem_bus_in_14( io_mem_bus_in_14 ),
       .io_mem_bus_in_13( io_mem_bus_in_13 ),
       .io_mem_bus_in_12( io_mem_bus_in_12 ),
       .io_mem_bus_in_11( io_mem_bus_in_11 ),
       .io_mem_bus_in_10( io_mem_bus_in_10 ),
       .io_mem_bus_in_9( io_mem_bus_in_9 ),
       .io_mem_bus_in_8( io_mem_bus_in_8 ),
       .io_mem_bus_in_7( io_mem_bus_in_7 ),
       .io_mem_bus_in_6( io_mem_bus_in_6 ),
       .io_mem_bus_in_5( io_mem_bus_in_5 ),
       .io_mem_bus_in_4( io_mem_bus_in_4 ),
       .io_mem_bus_in_3( io_mem_bus_in_3 ),
       .io_mem_bus_in_2( io_mem_bus_in_2 ),
       .io_mem_bus_in_1( io_mem_bus_in_1 ),
       .io_mem_bus_in_0( io_mem_bus_in_0 ),
       .io_H_out_above_22( T1498 ),
       .io_H_out_above_21( T1497 ),
       .io_H_out_above_20( T1496 ),
       .io_H_out_above_19( T1495 ),
       .io_H_out_above_18( T1494 ),
       .io_H_out_above_17( T1493 ),
       .io_H_out_above_16( T1492 ),
       .io_H_out_above_15( T1491 ),
       .io_H_out_above_14( T1490 ),
       .io_H_out_above_13( T1489 ),
       .io_H_out_above_12( T1488 ),
       .io_H_out_above_11( T1487 ),
       .io_H_out_above_10( T1486 ),
       .io_H_out_above_9( T1485 ),
       .io_H_out_above_8( T1484 ),
       .io_H_out_above_7( T1483 ),
       .io_H_out_above_6( T1482 ),
       .io_H_out_above_5( T1481 ),
       .io_H_out_above_4( T1480 ),
       .io_H_out_above_3( T1479 ),
       .io_H_out_above_2( T1478 ),
       .io_H_out_above_1( T1477 ),
       .io_H_out_above_0( T1476 ),
       .io_H_out_22( ArrayRowModule_io_H_out_22 ),
       .io_H_out_21( ArrayRowModule_io_H_out_21 ),
       .io_H_out_20( ArrayRowModule_io_H_out_20 ),
       .io_H_out_19( ArrayRowModule_io_H_out_19 ),
       .io_H_out_18( ArrayRowModule_io_H_out_18 ),
       .io_H_out_17( ArrayRowModule_io_H_out_17 ),
       .io_H_out_16( ArrayRowModule_io_H_out_16 ),
       .io_H_out_15( ArrayRowModule_io_H_out_15 ),
       .io_H_out_14( ArrayRowModule_io_H_out_14 ),
       .io_H_out_13( ArrayRowModule_io_H_out_13 ),
       .io_H_out_12( ArrayRowModule_io_H_out_12 ),
       .io_H_out_11( ArrayRowModule_io_H_out_11 ),
       .io_H_out_10( ArrayRowModule_io_H_out_10 ),
       .io_H_out_9( ArrayRowModule_io_H_out_9 ),
       .io_H_out_8( ArrayRowModule_io_H_out_8 ),
       .io_H_out_7( ArrayRowModule_io_H_out_7 ),
       .io_H_out_6( ArrayRowModule_io_H_out_6 ),
       .io_H_out_5( ArrayRowModule_io_H_out_5 ),
       .io_H_out_4( ArrayRowModule_io_H_out_4 ),
       .io_H_out_3( ArrayRowModule_io_H_out_3 ),
       .io_H_out_2( ArrayRowModule_io_H_out_2 ),
       .io_H_out_1( ArrayRowModule_io_H_out_1 ),
       .io_H_out_0( ArrayRowModule_io_H_out_0 ),
       .io_G_wire_below_3( ArrayRowModule_io_G_wire_below_3 ),
       .io_G_wire_below_2( ArrayRowModule_io_G_wire_below_2 ),
       .io_G_wire_below_1( ArrayRowModule_io_G_wire_below_1 ),
       .io_G_wire_below_0( ArrayRowModule_io_G_wire_below_0 ),
       .io_H_wire_below_32( ArrayRowModule_io_H_wire_below_32 ),
       .io_H_wire_below_31( ArrayRowModule_io_H_wire_below_31 ),
       .io_H_wire_below_30( ArrayRowModule_io_H_wire_below_30 ),
       .io_H_wire_below_29( ArrayRowModule_io_H_wire_below_29 ),
       .io_H_wire_below_28( ArrayRowModule_io_H_wire_below_28 ),
       .io_H_wire_below_27( ArrayRowModule_io_H_wire_below_27 ),
       .io_H_wire_below_26( ArrayRowModule_io_H_wire_below_26 ),
       .io_H_wire_below_25( ArrayRowModule_io_H_wire_below_25 ),
       .io_H_wire_below_24( ArrayRowModule_io_H_wire_below_24 ),
       .io_H_wire_below_23( ArrayRowModule_io_H_wire_below_23 ),
       .io_H_wire_below_22( ArrayRowModule_io_H_wire_below_22 ),
       .io_H_wire_below_21( ArrayRowModule_io_H_wire_below_21 ),
       .io_H_wire_below_20( ArrayRowModule_io_H_wire_below_20 ),
       .io_H_wire_below_19( ArrayRowModule_io_H_wire_below_19 ),
       .io_H_wire_below_18( ArrayRowModule_io_H_wire_below_18 ),
       .io_H_wire_below_17( ArrayRowModule_io_H_wire_below_17 ),
       .io_H_wire_below_16( ArrayRowModule_io_H_wire_below_16 ),
       .io_H_wire_below_15( ArrayRowModule_io_H_wire_below_15 ),
       .io_H_wire_below_14( ArrayRowModule_io_H_wire_below_14 ),
       .io_H_wire_below_13( ArrayRowModule_io_H_wire_below_13 ),
       .io_H_wire_below_12( ArrayRowModule_io_H_wire_below_12 ),
       .io_H_wire_below_11( ArrayRowModule_io_H_wire_below_11 ),
       .io_H_wire_below_10( ArrayRowModule_io_H_wire_below_10 ),
       .io_H_wire_below_9( ArrayRowModule_io_H_wire_below_9 ),
       .io_H_wire_below_8( ArrayRowModule_io_H_wire_below_8 ),
       .io_H_wire_below_7( ArrayRowModule_io_H_wire_below_7 ),
       .io_H_wire_below_6( ArrayRowModule_io_H_wire_below_6 ),
       .io_H_wire_below_5( ArrayRowModule_io_H_wire_below_5 ),
       .io_H_wire_below_4( ArrayRowModule_io_H_wire_below_4 ),
       .io_H_wire_below_3( ArrayRowModule_io_H_wire_below_3 ),
       .io_H_wire_below_2( ArrayRowModule_io_H_wire_below_2 ),
       .io_H_wire_below_1( ArrayRowModule_io_H_wire_below_1 ),
       .io_H_wire_below_0( ArrayRowModule_io_H_wire_below_0 ),
       .io_row_en( T1475 ),
       //.io_config_or_load(  )
       //.io_D_or_Z(  )
       .io_mem_bus_out_23( ArrayRowModule_io_mem_bus_out_23 ),
       .io_mem_bus_out_22( ArrayRowModule_io_mem_bus_out_22 ),
       .io_mem_bus_out_21( ArrayRowModule_io_mem_bus_out_21 ),
       .io_mem_bus_out_20( ArrayRowModule_io_mem_bus_out_20 ),
       .io_mem_bus_out_19( ArrayRowModule_io_mem_bus_out_19 ),
       .io_mem_bus_out_18( ArrayRowModule_io_mem_bus_out_18 ),
       .io_mem_bus_out_17( ArrayRowModule_io_mem_bus_out_17 ),
       .io_mem_bus_out_16( ArrayRowModule_io_mem_bus_out_16 ),
       .io_mem_bus_out_15( ArrayRowModule_io_mem_bus_out_15 ),
       .io_mem_bus_out_14( ArrayRowModule_io_mem_bus_out_14 ),
       .io_mem_bus_out_13( ArrayRowModule_io_mem_bus_out_13 ),
       .io_mem_bus_out_12( ArrayRowModule_io_mem_bus_out_12 ),
       .io_mem_bus_out_11( ArrayRowModule_io_mem_bus_out_11 ),
       .io_mem_bus_out_10( ArrayRowModule_io_mem_bus_out_10 ),
       .io_mem_bus_out_9( ArrayRowModule_io_mem_bus_out_9 ),
       .io_mem_bus_out_8( ArrayRowModule_io_mem_bus_out_8 ),
       .io_mem_bus_out_7( ArrayRowModule_io_mem_bus_out_7 ),
       .io_mem_bus_out_6( ArrayRowModule_io_mem_bus_out_6 ),
       .io_mem_bus_out_5( ArrayRowModule_io_mem_bus_out_5 ),
       .io_mem_bus_out_4( ArrayRowModule_io_mem_bus_out_4 ),
       .io_mem_bus_out_3( ArrayRowModule_io_mem_bus_out_3 ),
       .io_mem_bus_out_2( ArrayRowModule_io_mem_bus_out_2 ),
       .io_mem_bus_out_1( ArrayRowModule_io_mem_bus_out_1 ),
       .io_mem_bus_out_0( ArrayRowModule_io_mem_bus_out_0 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ArrayRowModule.io_config_or_load = {1{$random}};
    assign ArrayRowModule.io_D_or_Z = {1{$random}};
    assign ArrayRowModule.io_mem_bus_out_23 = {1{$random}};
// synthesis translate_on
`endif
  ArrayRowModule ArrayRowModule_1(.clk(clk), .reset(reset),
       .io_V_wire_in_367( VwireModule_io_VwirePorts_1_22_15_out ),
       .io_V_wire_in_366( VwireModule_io_VwirePorts_1_22_14_out ),
       .io_V_wire_in_365( VwireModule_io_VwirePorts_1_22_13_out ),
       .io_V_wire_in_364( VwireModule_io_VwirePorts_1_22_12_out ),
       .io_V_wire_in_363( VwireModule_io_VwirePorts_1_22_11_out ),
       .io_V_wire_in_362( VwireModule_io_VwirePorts_1_22_10_out ),
       .io_V_wire_in_361( VwireModule_io_VwirePorts_1_22_9_out ),
       .io_V_wire_in_360( VwireModule_io_VwirePorts_1_22_8_out ),
       .io_V_wire_in_359( VwireModule_io_VwirePorts_1_22_7_out ),
       .io_V_wire_in_358( VwireModule_io_VwirePorts_1_22_6_out ),
       .io_V_wire_in_357( VwireModule_io_VwirePorts_1_22_5_out ),
       .io_V_wire_in_356( VwireModule_io_VwirePorts_1_22_4_out ),
       .io_V_wire_in_355( VwireModule_io_VwirePorts_1_22_3_out ),
       .io_V_wire_in_354( VwireModule_io_VwirePorts_1_22_2_out ),
       .io_V_wire_in_353( VwireModule_io_VwirePorts_1_22_1_out ),
       .io_V_wire_in_352( VwireModule_io_VwirePorts_1_22_0_out ),
       .io_V_wire_in_351( VwireModule_io_VwirePorts_1_21_15_out ),
       .io_V_wire_in_350( VwireModule_io_VwirePorts_1_21_14_out ),
       .io_V_wire_in_349( VwireModule_io_VwirePorts_1_21_13_out ),
       .io_V_wire_in_348( VwireModule_io_VwirePorts_1_21_12_out ),
       .io_V_wire_in_347( VwireModule_io_VwirePorts_1_21_11_out ),
       .io_V_wire_in_346( VwireModule_io_VwirePorts_1_21_10_out ),
       .io_V_wire_in_345( VwireModule_io_VwirePorts_1_21_9_out ),
       .io_V_wire_in_344( VwireModule_io_VwirePorts_1_21_8_out ),
       .io_V_wire_in_343( VwireModule_io_VwirePorts_1_21_7_out ),
       .io_V_wire_in_342( VwireModule_io_VwirePorts_1_21_6_out ),
       .io_V_wire_in_341( VwireModule_io_VwirePorts_1_21_5_out ),
       .io_V_wire_in_340( VwireModule_io_VwirePorts_1_21_4_out ),
       .io_V_wire_in_339( VwireModule_io_VwirePorts_1_21_3_out ),
       .io_V_wire_in_338( VwireModule_io_VwirePorts_1_21_2_out ),
       .io_V_wire_in_337( VwireModule_io_VwirePorts_1_21_1_out ),
       .io_V_wire_in_336( VwireModule_io_VwirePorts_1_21_0_out ),
       .io_V_wire_in_335( VwireModule_io_VwirePorts_1_20_15_out ),
       .io_V_wire_in_334( VwireModule_io_VwirePorts_1_20_14_out ),
       .io_V_wire_in_333( VwireModule_io_VwirePorts_1_20_13_out ),
       .io_V_wire_in_332( VwireModule_io_VwirePorts_1_20_12_out ),
       .io_V_wire_in_331( VwireModule_io_VwirePorts_1_20_11_out ),
       .io_V_wire_in_330( VwireModule_io_VwirePorts_1_20_10_out ),
       .io_V_wire_in_329( VwireModule_io_VwirePorts_1_20_9_out ),
       .io_V_wire_in_328( VwireModule_io_VwirePorts_1_20_8_out ),
       .io_V_wire_in_327( VwireModule_io_VwirePorts_1_20_7_out ),
       .io_V_wire_in_326( VwireModule_io_VwirePorts_1_20_6_out ),
       .io_V_wire_in_325( VwireModule_io_VwirePorts_1_20_5_out ),
       .io_V_wire_in_324( VwireModule_io_VwirePorts_1_20_4_out ),
       .io_V_wire_in_323( VwireModule_io_VwirePorts_1_20_3_out ),
       .io_V_wire_in_322( VwireModule_io_VwirePorts_1_20_2_out ),
       .io_V_wire_in_321( VwireModule_io_VwirePorts_1_20_1_out ),
       .io_V_wire_in_320( VwireModule_io_VwirePorts_1_20_0_out ),
       .io_V_wire_in_319( VwireModule_io_VwirePorts_1_19_15_out ),
       .io_V_wire_in_318( VwireModule_io_VwirePorts_1_19_14_out ),
       .io_V_wire_in_317( VwireModule_io_VwirePorts_1_19_13_out ),
       .io_V_wire_in_316( VwireModule_io_VwirePorts_1_19_12_out ),
       .io_V_wire_in_315( VwireModule_io_VwirePorts_1_19_11_out ),
       .io_V_wire_in_314( VwireModule_io_VwirePorts_1_19_10_out ),
       .io_V_wire_in_313( VwireModule_io_VwirePorts_1_19_9_out ),
       .io_V_wire_in_312( VwireModule_io_VwirePorts_1_19_8_out ),
       .io_V_wire_in_311( VwireModule_io_VwirePorts_1_19_7_out ),
       .io_V_wire_in_310( VwireModule_io_VwirePorts_1_19_6_out ),
       .io_V_wire_in_309( VwireModule_io_VwirePorts_1_19_5_out ),
       .io_V_wire_in_308( VwireModule_io_VwirePorts_1_19_4_out ),
       .io_V_wire_in_307( VwireModule_io_VwirePorts_1_19_3_out ),
       .io_V_wire_in_306( VwireModule_io_VwirePorts_1_19_2_out ),
       .io_V_wire_in_305( VwireModule_io_VwirePorts_1_19_1_out ),
       .io_V_wire_in_304( VwireModule_io_VwirePorts_1_19_0_out ),
       .io_V_wire_in_303( VwireModule_io_VwirePorts_1_18_15_out ),
       .io_V_wire_in_302( VwireModule_io_VwirePorts_1_18_14_out ),
       .io_V_wire_in_301( VwireModule_io_VwirePorts_1_18_13_out ),
       .io_V_wire_in_300( VwireModule_io_VwirePorts_1_18_12_out ),
       .io_V_wire_in_299( VwireModule_io_VwirePorts_1_18_11_out ),
       .io_V_wire_in_298( VwireModule_io_VwirePorts_1_18_10_out ),
       .io_V_wire_in_297( VwireModule_io_VwirePorts_1_18_9_out ),
       .io_V_wire_in_296( VwireModule_io_VwirePorts_1_18_8_out ),
       .io_V_wire_in_295( VwireModule_io_VwirePorts_1_18_7_out ),
       .io_V_wire_in_294( VwireModule_io_VwirePorts_1_18_6_out ),
       .io_V_wire_in_293( VwireModule_io_VwirePorts_1_18_5_out ),
       .io_V_wire_in_292( VwireModule_io_VwirePorts_1_18_4_out ),
       .io_V_wire_in_291( VwireModule_io_VwirePorts_1_18_3_out ),
       .io_V_wire_in_290( VwireModule_io_VwirePorts_1_18_2_out ),
       .io_V_wire_in_289( VwireModule_io_VwirePorts_1_18_1_out ),
       .io_V_wire_in_288( VwireModule_io_VwirePorts_1_18_0_out ),
       .io_V_wire_in_287( VwireModule_io_VwirePorts_1_17_15_out ),
       .io_V_wire_in_286( VwireModule_io_VwirePorts_1_17_14_out ),
       .io_V_wire_in_285( VwireModule_io_VwirePorts_1_17_13_out ),
       .io_V_wire_in_284( VwireModule_io_VwirePorts_1_17_12_out ),
       .io_V_wire_in_283( VwireModule_io_VwirePorts_1_17_11_out ),
       .io_V_wire_in_282( VwireModule_io_VwirePorts_1_17_10_out ),
       .io_V_wire_in_281( VwireModule_io_VwirePorts_1_17_9_out ),
       .io_V_wire_in_280( VwireModule_io_VwirePorts_1_17_8_out ),
       .io_V_wire_in_279( VwireModule_io_VwirePorts_1_17_7_out ),
       .io_V_wire_in_278( VwireModule_io_VwirePorts_1_17_6_out ),
       .io_V_wire_in_277( VwireModule_io_VwirePorts_1_17_5_out ),
       .io_V_wire_in_276( VwireModule_io_VwirePorts_1_17_4_out ),
       .io_V_wire_in_275( VwireModule_io_VwirePorts_1_17_3_out ),
       .io_V_wire_in_274( VwireModule_io_VwirePorts_1_17_2_out ),
       .io_V_wire_in_273( VwireModule_io_VwirePorts_1_17_1_out ),
       .io_V_wire_in_272( VwireModule_io_VwirePorts_1_17_0_out ),
       .io_V_wire_in_271( VwireModule_io_VwirePorts_1_16_15_out ),
       .io_V_wire_in_270( VwireModule_io_VwirePorts_1_16_14_out ),
       .io_V_wire_in_269( VwireModule_io_VwirePorts_1_16_13_out ),
       .io_V_wire_in_268( VwireModule_io_VwirePorts_1_16_12_out ),
       .io_V_wire_in_267( VwireModule_io_VwirePorts_1_16_11_out ),
       .io_V_wire_in_266( VwireModule_io_VwirePorts_1_16_10_out ),
       .io_V_wire_in_265( VwireModule_io_VwirePorts_1_16_9_out ),
       .io_V_wire_in_264( VwireModule_io_VwirePorts_1_16_8_out ),
       .io_V_wire_in_263( VwireModule_io_VwirePorts_1_16_7_out ),
       .io_V_wire_in_262( VwireModule_io_VwirePorts_1_16_6_out ),
       .io_V_wire_in_261( VwireModule_io_VwirePorts_1_16_5_out ),
       .io_V_wire_in_260( VwireModule_io_VwirePorts_1_16_4_out ),
       .io_V_wire_in_259( VwireModule_io_VwirePorts_1_16_3_out ),
       .io_V_wire_in_258( VwireModule_io_VwirePorts_1_16_2_out ),
       .io_V_wire_in_257( VwireModule_io_VwirePorts_1_16_1_out ),
       .io_V_wire_in_256( VwireModule_io_VwirePorts_1_16_0_out ),
       .io_V_wire_in_255( VwireModule_io_VwirePorts_1_15_15_out ),
       .io_V_wire_in_254( VwireModule_io_VwirePorts_1_15_14_out ),
       .io_V_wire_in_253( VwireModule_io_VwirePorts_1_15_13_out ),
       .io_V_wire_in_252( VwireModule_io_VwirePorts_1_15_12_out ),
       .io_V_wire_in_251( VwireModule_io_VwirePorts_1_15_11_out ),
       .io_V_wire_in_250( VwireModule_io_VwirePorts_1_15_10_out ),
       .io_V_wire_in_249( VwireModule_io_VwirePorts_1_15_9_out ),
       .io_V_wire_in_248( VwireModule_io_VwirePorts_1_15_8_out ),
       .io_V_wire_in_247( VwireModule_io_VwirePorts_1_15_7_out ),
       .io_V_wire_in_246( VwireModule_io_VwirePorts_1_15_6_out ),
       .io_V_wire_in_245( VwireModule_io_VwirePorts_1_15_5_out ),
       .io_V_wire_in_244( VwireModule_io_VwirePorts_1_15_4_out ),
       .io_V_wire_in_243( VwireModule_io_VwirePorts_1_15_3_out ),
       .io_V_wire_in_242( VwireModule_io_VwirePorts_1_15_2_out ),
       .io_V_wire_in_241( VwireModule_io_VwirePorts_1_15_1_out ),
       .io_V_wire_in_240( VwireModule_io_VwirePorts_1_15_0_out ),
       .io_V_wire_in_239( VwireModule_io_VwirePorts_1_14_15_out ),
       .io_V_wire_in_238( VwireModule_io_VwirePorts_1_14_14_out ),
       .io_V_wire_in_237( VwireModule_io_VwirePorts_1_14_13_out ),
       .io_V_wire_in_236( VwireModule_io_VwirePorts_1_14_12_out ),
       .io_V_wire_in_235( VwireModule_io_VwirePorts_1_14_11_out ),
       .io_V_wire_in_234( VwireModule_io_VwirePorts_1_14_10_out ),
       .io_V_wire_in_233( VwireModule_io_VwirePorts_1_14_9_out ),
       .io_V_wire_in_232( VwireModule_io_VwirePorts_1_14_8_out ),
       .io_V_wire_in_231( VwireModule_io_VwirePorts_1_14_7_out ),
       .io_V_wire_in_230( VwireModule_io_VwirePorts_1_14_6_out ),
       .io_V_wire_in_229( VwireModule_io_VwirePorts_1_14_5_out ),
       .io_V_wire_in_228( VwireModule_io_VwirePorts_1_14_4_out ),
       .io_V_wire_in_227( VwireModule_io_VwirePorts_1_14_3_out ),
       .io_V_wire_in_226( VwireModule_io_VwirePorts_1_14_2_out ),
       .io_V_wire_in_225( VwireModule_io_VwirePorts_1_14_1_out ),
       .io_V_wire_in_224( VwireModule_io_VwirePorts_1_14_0_out ),
       .io_V_wire_in_223( VwireModule_io_VwirePorts_1_13_15_out ),
       .io_V_wire_in_222( VwireModule_io_VwirePorts_1_13_14_out ),
       .io_V_wire_in_221( VwireModule_io_VwirePorts_1_13_13_out ),
       .io_V_wire_in_220( VwireModule_io_VwirePorts_1_13_12_out ),
       .io_V_wire_in_219( VwireModule_io_VwirePorts_1_13_11_out ),
       .io_V_wire_in_218( VwireModule_io_VwirePorts_1_13_10_out ),
       .io_V_wire_in_217( VwireModule_io_VwirePorts_1_13_9_out ),
       .io_V_wire_in_216( VwireModule_io_VwirePorts_1_13_8_out ),
       .io_V_wire_in_215( VwireModule_io_VwirePorts_1_13_7_out ),
       .io_V_wire_in_214( VwireModule_io_VwirePorts_1_13_6_out ),
       .io_V_wire_in_213( VwireModule_io_VwirePorts_1_13_5_out ),
       .io_V_wire_in_212( VwireModule_io_VwirePorts_1_13_4_out ),
       .io_V_wire_in_211( VwireModule_io_VwirePorts_1_13_3_out ),
       .io_V_wire_in_210( VwireModule_io_VwirePorts_1_13_2_out ),
       .io_V_wire_in_209( VwireModule_io_VwirePorts_1_13_1_out ),
       .io_V_wire_in_208( VwireModule_io_VwirePorts_1_13_0_out ),
       .io_V_wire_in_207( VwireModule_io_VwirePorts_1_12_15_out ),
       .io_V_wire_in_206( VwireModule_io_VwirePorts_1_12_14_out ),
       .io_V_wire_in_205( VwireModule_io_VwirePorts_1_12_13_out ),
       .io_V_wire_in_204( VwireModule_io_VwirePorts_1_12_12_out ),
       .io_V_wire_in_203( VwireModule_io_VwirePorts_1_12_11_out ),
       .io_V_wire_in_202( VwireModule_io_VwirePorts_1_12_10_out ),
       .io_V_wire_in_201( VwireModule_io_VwirePorts_1_12_9_out ),
       .io_V_wire_in_200( VwireModule_io_VwirePorts_1_12_8_out ),
       .io_V_wire_in_199( VwireModule_io_VwirePorts_1_12_7_out ),
       .io_V_wire_in_198( VwireModule_io_VwirePorts_1_12_6_out ),
       .io_V_wire_in_197( VwireModule_io_VwirePorts_1_12_5_out ),
       .io_V_wire_in_196( VwireModule_io_VwirePorts_1_12_4_out ),
       .io_V_wire_in_195( VwireModule_io_VwirePorts_1_12_3_out ),
       .io_V_wire_in_194( VwireModule_io_VwirePorts_1_12_2_out ),
       .io_V_wire_in_193( VwireModule_io_VwirePorts_1_12_1_out ),
       .io_V_wire_in_192( VwireModule_io_VwirePorts_1_12_0_out ),
       .io_V_wire_in_191( VwireModule_io_VwirePorts_1_11_15_out ),
       .io_V_wire_in_190( VwireModule_io_VwirePorts_1_11_14_out ),
       .io_V_wire_in_189( VwireModule_io_VwirePorts_1_11_13_out ),
       .io_V_wire_in_188( VwireModule_io_VwirePorts_1_11_12_out ),
       .io_V_wire_in_187( VwireModule_io_VwirePorts_1_11_11_out ),
       .io_V_wire_in_186( VwireModule_io_VwirePorts_1_11_10_out ),
       .io_V_wire_in_185( VwireModule_io_VwirePorts_1_11_9_out ),
       .io_V_wire_in_184( VwireModule_io_VwirePorts_1_11_8_out ),
       .io_V_wire_in_183( VwireModule_io_VwirePorts_1_11_7_out ),
       .io_V_wire_in_182( VwireModule_io_VwirePorts_1_11_6_out ),
       .io_V_wire_in_181( VwireModule_io_VwirePorts_1_11_5_out ),
       .io_V_wire_in_180( VwireModule_io_VwirePorts_1_11_4_out ),
       .io_V_wire_in_179( VwireModule_io_VwirePorts_1_11_3_out ),
       .io_V_wire_in_178( VwireModule_io_VwirePorts_1_11_2_out ),
       .io_V_wire_in_177( VwireModule_io_VwirePorts_1_11_1_out ),
       .io_V_wire_in_176( VwireModule_io_VwirePorts_1_11_0_out ),
       .io_V_wire_in_175( VwireModule_io_VwirePorts_1_10_15_out ),
       .io_V_wire_in_174( VwireModule_io_VwirePorts_1_10_14_out ),
       .io_V_wire_in_173( VwireModule_io_VwirePorts_1_10_13_out ),
       .io_V_wire_in_172( VwireModule_io_VwirePorts_1_10_12_out ),
       .io_V_wire_in_171( VwireModule_io_VwirePorts_1_10_11_out ),
       .io_V_wire_in_170( VwireModule_io_VwirePorts_1_10_10_out ),
       .io_V_wire_in_169( VwireModule_io_VwirePorts_1_10_9_out ),
       .io_V_wire_in_168( VwireModule_io_VwirePorts_1_10_8_out ),
       .io_V_wire_in_167( VwireModule_io_VwirePorts_1_10_7_out ),
       .io_V_wire_in_166( VwireModule_io_VwirePorts_1_10_6_out ),
       .io_V_wire_in_165( VwireModule_io_VwirePorts_1_10_5_out ),
       .io_V_wire_in_164( VwireModule_io_VwirePorts_1_10_4_out ),
       .io_V_wire_in_163( VwireModule_io_VwirePorts_1_10_3_out ),
       .io_V_wire_in_162( VwireModule_io_VwirePorts_1_10_2_out ),
       .io_V_wire_in_161( VwireModule_io_VwirePorts_1_10_1_out ),
       .io_V_wire_in_160( VwireModule_io_VwirePorts_1_10_0_out ),
       .io_V_wire_in_159( VwireModule_io_VwirePorts_1_9_15_out ),
       .io_V_wire_in_158( VwireModule_io_VwirePorts_1_9_14_out ),
       .io_V_wire_in_157( VwireModule_io_VwirePorts_1_9_13_out ),
       .io_V_wire_in_156( VwireModule_io_VwirePorts_1_9_12_out ),
       .io_V_wire_in_155( VwireModule_io_VwirePorts_1_9_11_out ),
       .io_V_wire_in_154( VwireModule_io_VwirePorts_1_9_10_out ),
       .io_V_wire_in_153( VwireModule_io_VwirePorts_1_9_9_out ),
       .io_V_wire_in_152( VwireModule_io_VwirePorts_1_9_8_out ),
       .io_V_wire_in_151( VwireModule_io_VwirePorts_1_9_7_out ),
       .io_V_wire_in_150( VwireModule_io_VwirePorts_1_9_6_out ),
       .io_V_wire_in_149( VwireModule_io_VwirePorts_1_9_5_out ),
       .io_V_wire_in_148( VwireModule_io_VwirePorts_1_9_4_out ),
       .io_V_wire_in_147( VwireModule_io_VwirePorts_1_9_3_out ),
       .io_V_wire_in_146( VwireModule_io_VwirePorts_1_9_2_out ),
       .io_V_wire_in_145( VwireModule_io_VwirePorts_1_9_1_out ),
       .io_V_wire_in_144( VwireModule_io_VwirePorts_1_9_0_out ),
       .io_V_wire_in_143( VwireModule_io_VwirePorts_1_8_15_out ),
       .io_V_wire_in_142( VwireModule_io_VwirePorts_1_8_14_out ),
       .io_V_wire_in_141( VwireModule_io_VwirePorts_1_8_13_out ),
       .io_V_wire_in_140( VwireModule_io_VwirePorts_1_8_12_out ),
       .io_V_wire_in_139( VwireModule_io_VwirePorts_1_8_11_out ),
       .io_V_wire_in_138( VwireModule_io_VwirePorts_1_8_10_out ),
       .io_V_wire_in_137( VwireModule_io_VwirePorts_1_8_9_out ),
       .io_V_wire_in_136( VwireModule_io_VwirePorts_1_8_8_out ),
       .io_V_wire_in_135( VwireModule_io_VwirePorts_1_8_7_out ),
       .io_V_wire_in_134( VwireModule_io_VwirePorts_1_8_6_out ),
       .io_V_wire_in_133( VwireModule_io_VwirePorts_1_8_5_out ),
       .io_V_wire_in_132( VwireModule_io_VwirePorts_1_8_4_out ),
       .io_V_wire_in_131( VwireModule_io_VwirePorts_1_8_3_out ),
       .io_V_wire_in_130( VwireModule_io_VwirePorts_1_8_2_out ),
       .io_V_wire_in_129( VwireModule_io_VwirePorts_1_8_1_out ),
       .io_V_wire_in_128( VwireModule_io_VwirePorts_1_8_0_out ),
       .io_V_wire_in_127( VwireModule_io_VwirePorts_1_7_15_out ),
       .io_V_wire_in_126( VwireModule_io_VwirePorts_1_7_14_out ),
       .io_V_wire_in_125( VwireModule_io_VwirePorts_1_7_13_out ),
       .io_V_wire_in_124( VwireModule_io_VwirePorts_1_7_12_out ),
       .io_V_wire_in_123( VwireModule_io_VwirePorts_1_7_11_out ),
       .io_V_wire_in_122( VwireModule_io_VwirePorts_1_7_10_out ),
       .io_V_wire_in_121( VwireModule_io_VwirePorts_1_7_9_out ),
       .io_V_wire_in_120( VwireModule_io_VwirePorts_1_7_8_out ),
       .io_V_wire_in_119( VwireModule_io_VwirePorts_1_7_7_out ),
       .io_V_wire_in_118( VwireModule_io_VwirePorts_1_7_6_out ),
       .io_V_wire_in_117( VwireModule_io_VwirePorts_1_7_5_out ),
       .io_V_wire_in_116( VwireModule_io_VwirePorts_1_7_4_out ),
       .io_V_wire_in_115( VwireModule_io_VwirePorts_1_7_3_out ),
       .io_V_wire_in_114( VwireModule_io_VwirePorts_1_7_2_out ),
       .io_V_wire_in_113( VwireModule_io_VwirePorts_1_7_1_out ),
       .io_V_wire_in_112( VwireModule_io_VwirePorts_1_7_0_out ),
       .io_V_wire_in_111( VwireModule_io_VwirePorts_1_6_15_out ),
       .io_V_wire_in_110( VwireModule_io_VwirePorts_1_6_14_out ),
       .io_V_wire_in_109( VwireModule_io_VwirePorts_1_6_13_out ),
       .io_V_wire_in_108( VwireModule_io_VwirePorts_1_6_12_out ),
       .io_V_wire_in_107( VwireModule_io_VwirePorts_1_6_11_out ),
       .io_V_wire_in_106( VwireModule_io_VwirePorts_1_6_10_out ),
       .io_V_wire_in_105( VwireModule_io_VwirePorts_1_6_9_out ),
       .io_V_wire_in_104( VwireModule_io_VwirePorts_1_6_8_out ),
       .io_V_wire_in_103( VwireModule_io_VwirePorts_1_6_7_out ),
       .io_V_wire_in_102( VwireModule_io_VwirePorts_1_6_6_out ),
       .io_V_wire_in_101( VwireModule_io_VwirePorts_1_6_5_out ),
       .io_V_wire_in_100( VwireModule_io_VwirePorts_1_6_4_out ),
       .io_V_wire_in_99( VwireModule_io_VwirePorts_1_6_3_out ),
       .io_V_wire_in_98( VwireModule_io_VwirePorts_1_6_2_out ),
       .io_V_wire_in_97( VwireModule_io_VwirePorts_1_6_1_out ),
       .io_V_wire_in_96( VwireModule_io_VwirePorts_1_6_0_out ),
       .io_V_wire_in_95( VwireModule_io_VwirePorts_1_5_15_out ),
       .io_V_wire_in_94( VwireModule_io_VwirePorts_1_5_14_out ),
       .io_V_wire_in_93( VwireModule_io_VwirePorts_1_5_13_out ),
       .io_V_wire_in_92( VwireModule_io_VwirePorts_1_5_12_out ),
       .io_V_wire_in_91( VwireModule_io_VwirePorts_1_5_11_out ),
       .io_V_wire_in_90( VwireModule_io_VwirePorts_1_5_10_out ),
       .io_V_wire_in_89( VwireModule_io_VwirePorts_1_5_9_out ),
       .io_V_wire_in_88( VwireModule_io_VwirePorts_1_5_8_out ),
       .io_V_wire_in_87( VwireModule_io_VwirePorts_1_5_7_out ),
       .io_V_wire_in_86( VwireModule_io_VwirePorts_1_5_6_out ),
       .io_V_wire_in_85( VwireModule_io_VwirePorts_1_5_5_out ),
       .io_V_wire_in_84( VwireModule_io_VwirePorts_1_5_4_out ),
       .io_V_wire_in_83( VwireModule_io_VwirePorts_1_5_3_out ),
       .io_V_wire_in_82( VwireModule_io_VwirePorts_1_5_2_out ),
       .io_V_wire_in_81( VwireModule_io_VwirePorts_1_5_1_out ),
       .io_V_wire_in_80( VwireModule_io_VwirePorts_1_5_0_out ),
       .io_V_wire_in_79( VwireModule_io_VwirePorts_1_4_15_out ),
       .io_V_wire_in_78( VwireModule_io_VwirePorts_1_4_14_out ),
       .io_V_wire_in_77( VwireModule_io_VwirePorts_1_4_13_out ),
       .io_V_wire_in_76( VwireModule_io_VwirePorts_1_4_12_out ),
       .io_V_wire_in_75( VwireModule_io_VwirePorts_1_4_11_out ),
       .io_V_wire_in_74( VwireModule_io_VwirePorts_1_4_10_out ),
       .io_V_wire_in_73( VwireModule_io_VwirePorts_1_4_9_out ),
       .io_V_wire_in_72( VwireModule_io_VwirePorts_1_4_8_out ),
       .io_V_wire_in_71( VwireModule_io_VwirePorts_1_4_7_out ),
       .io_V_wire_in_70( VwireModule_io_VwirePorts_1_4_6_out ),
       .io_V_wire_in_69( VwireModule_io_VwirePorts_1_4_5_out ),
       .io_V_wire_in_68( VwireModule_io_VwirePorts_1_4_4_out ),
       .io_V_wire_in_67( VwireModule_io_VwirePorts_1_4_3_out ),
       .io_V_wire_in_66( VwireModule_io_VwirePorts_1_4_2_out ),
       .io_V_wire_in_65( VwireModule_io_VwirePorts_1_4_1_out ),
       .io_V_wire_in_64( VwireModule_io_VwirePorts_1_4_0_out ),
       .io_V_wire_in_63( VwireModule_io_VwirePorts_1_3_15_out ),
       .io_V_wire_in_62( VwireModule_io_VwirePorts_1_3_14_out ),
       .io_V_wire_in_61( VwireModule_io_VwirePorts_1_3_13_out ),
       .io_V_wire_in_60( VwireModule_io_VwirePorts_1_3_12_out ),
       .io_V_wire_in_59( VwireModule_io_VwirePorts_1_3_11_out ),
       .io_V_wire_in_58( VwireModule_io_VwirePorts_1_3_10_out ),
       .io_V_wire_in_57( VwireModule_io_VwirePorts_1_3_9_out ),
       .io_V_wire_in_56( VwireModule_io_VwirePorts_1_3_8_out ),
       .io_V_wire_in_55( VwireModule_io_VwirePorts_1_3_7_out ),
       .io_V_wire_in_54( VwireModule_io_VwirePorts_1_3_6_out ),
       .io_V_wire_in_53( VwireModule_io_VwirePorts_1_3_5_out ),
       .io_V_wire_in_52( VwireModule_io_VwirePorts_1_3_4_out ),
       .io_V_wire_in_51( VwireModule_io_VwirePorts_1_3_3_out ),
       .io_V_wire_in_50( VwireModule_io_VwirePorts_1_3_2_out ),
       .io_V_wire_in_49( VwireModule_io_VwirePorts_1_3_1_out ),
       .io_V_wire_in_48( VwireModule_io_VwirePorts_1_3_0_out ),
       .io_V_wire_in_47( VwireModule_io_VwirePorts_1_2_15_out ),
       .io_V_wire_in_46( VwireModule_io_VwirePorts_1_2_14_out ),
       .io_V_wire_in_45( VwireModule_io_VwirePorts_1_2_13_out ),
       .io_V_wire_in_44( VwireModule_io_VwirePorts_1_2_12_out ),
       .io_V_wire_in_43( VwireModule_io_VwirePorts_1_2_11_out ),
       .io_V_wire_in_42( VwireModule_io_VwirePorts_1_2_10_out ),
       .io_V_wire_in_41( VwireModule_io_VwirePorts_1_2_9_out ),
       .io_V_wire_in_40( VwireModule_io_VwirePorts_1_2_8_out ),
       .io_V_wire_in_39( VwireModule_io_VwirePorts_1_2_7_out ),
       .io_V_wire_in_38( VwireModule_io_VwirePorts_1_2_6_out ),
       .io_V_wire_in_37( VwireModule_io_VwirePorts_1_2_5_out ),
       .io_V_wire_in_36( VwireModule_io_VwirePorts_1_2_4_out ),
       .io_V_wire_in_35( VwireModule_io_VwirePorts_1_2_3_out ),
       .io_V_wire_in_34( VwireModule_io_VwirePorts_1_2_2_out ),
       .io_V_wire_in_33( VwireModule_io_VwirePorts_1_2_1_out ),
       .io_V_wire_in_32( VwireModule_io_VwirePorts_1_2_0_out ),
       .io_V_wire_in_31( VwireModule_io_VwirePorts_1_1_15_out ),
       .io_V_wire_in_30( VwireModule_io_VwirePorts_1_1_14_out ),
       .io_V_wire_in_29( VwireModule_io_VwirePorts_1_1_13_out ),
       .io_V_wire_in_28( VwireModule_io_VwirePorts_1_1_12_out ),
       .io_V_wire_in_27( VwireModule_io_VwirePorts_1_1_11_out ),
       .io_V_wire_in_26( VwireModule_io_VwirePorts_1_1_10_out ),
       .io_V_wire_in_25( VwireModule_io_VwirePorts_1_1_9_out ),
       .io_V_wire_in_24( VwireModule_io_VwirePorts_1_1_8_out ),
       .io_V_wire_in_23( VwireModule_io_VwirePorts_1_1_7_out ),
       .io_V_wire_in_22( VwireModule_io_VwirePorts_1_1_6_out ),
       .io_V_wire_in_21( VwireModule_io_VwirePorts_1_1_5_out ),
       .io_V_wire_in_20( VwireModule_io_VwirePorts_1_1_4_out ),
       .io_V_wire_in_19( VwireModule_io_VwirePorts_1_1_3_out ),
       .io_V_wire_in_18( VwireModule_io_VwirePorts_1_1_2_out ),
       .io_V_wire_in_17( VwireModule_io_VwirePorts_1_1_1_out ),
       .io_V_wire_in_16( VwireModule_io_VwirePorts_1_1_0_out ),
       .io_V_wire_in_15( VwireModule_io_VwirePorts_1_0_15_out ),
       .io_V_wire_in_14( VwireModule_io_VwirePorts_1_0_14_out ),
       .io_V_wire_in_13( VwireModule_io_VwirePorts_1_0_13_out ),
       .io_V_wire_in_12( VwireModule_io_VwirePorts_1_0_12_out ),
       .io_V_wire_in_11( VwireModule_io_VwirePorts_1_0_11_out ),
       .io_V_wire_in_10( VwireModule_io_VwirePorts_1_0_10_out ),
       .io_V_wire_in_9( VwireModule_io_VwirePorts_1_0_9_out ),
       .io_V_wire_in_8( VwireModule_io_VwirePorts_1_0_8_out ),
       .io_V_wire_in_7( VwireModule_io_VwirePorts_1_0_7_out ),
       .io_V_wire_in_6( VwireModule_io_VwirePorts_1_0_6_out ),
       .io_V_wire_in_5( VwireModule_io_VwirePorts_1_0_5_out ),
       .io_V_wire_in_4( VwireModule_io_VwirePorts_1_0_4_out ),
       .io_V_wire_in_3( VwireModule_io_VwirePorts_1_0_3_out ),
       .io_V_wire_in_2( VwireModule_io_VwirePorts_1_0_2_out ),
       .io_V_wire_in_1( VwireModule_io_VwirePorts_1_0_1_out ),
       .io_V_wire_in_0( VwireModule_io_VwirePorts_1_0_0_out ),
       .io_V_wire_out_367( ArrayRowModule_1_io_V_wire_out_367 ),
       .io_V_wire_out_366( ArrayRowModule_1_io_V_wire_out_366 ),
       .io_V_wire_out_365( ArrayRowModule_1_io_V_wire_out_365 ),
       .io_V_wire_out_364( ArrayRowModule_1_io_V_wire_out_364 ),
       .io_V_wire_out_363( ArrayRowModule_1_io_V_wire_out_363 ),
       .io_V_wire_out_362( ArrayRowModule_1_io_V_wire_out_362 ),
       .io_V_wire_out_361( ArrayRowModule_1_io_V_wire_out_361 ),
       .io_V_wire_out_360( ArrayRowModule_1_io_V_wire_out_360 ),
       .io_V_wire_out_359( ArrayRowModule_1_io_V_wire_out_359 ),
       .io_V_wire_out_358( ArrayRowModule_1_io_V_wire_out_358 ),
       .io_V_wire_out_357( ArrayRowModule_1_io_V_wire_out_357 ),
       .io_V_wire_out_356( ArrayRowModule_1_io_V_wire_out_356 ),
       .io_V_wire_out_355( ArrayRowModule_1_io_V_wire_out_355 ),
       .io_V_wire_out_354( ArrayRowModule_1_io_V_wire_out_354 ),
       .io_V_wire_out_353( ArrayRowModule_1_io_V_wire_out_353 ),
       .io_V_wire_out_352( ArrayRowModule_1_io_V_wire_out_352 ),
       .io_V_wire_out_351( ArrayRowModule_1_io_V_wire_out_351 ),
       .io_V_wire_out_350( ArrayRowModule_1_io_V_wire_out_350 ),
       .io_V_wire_out_349( ArrayRowModule_1_io_V_wire_out_349 ),
       .io_V_wire_out_348( ArrayRowModule_1_io_V_wire_out_348 ),
       .io_V_wire_out_347( ArrayRowModule_1_io_V_wire_out_347 ),
       .io_V_wire_out_346( ArrayRowModule_1_io_V_wire_out_346 ),
       .io_V_wire_out_345( ArrayRowModule_1_io_V_wire_out_345 ),
       .io_V_wire_out_344( ArrayRowModule_1_io_V_wire_out_344 ),
       .io_V_wire_out_343( ArrayRowModule_1_io_V_wire_out_343 ),
       .io_V_wire_out_342( ArrayRowModule_1_io_V_wire_out_342 ),
       .io_V_wire_out_341( ArrayRowModule_1_io_V_wire_out_341 ),
       .io_V_wire_out_340( ArrayRowModule_1_io_V_wire_out_340 ),
       .io_V_wire_out_339( ArrayRowModule_1_io_V_wire_out_339 ),
       .io_V_wire_out_338( ArrayRowModule_1_io_V_wire_out_338 ),
       .io_V_wire_out_337( ArrayRowModule_1_io_V_wire_out_337 ),
       .io_V_wire_out_336( ArrayRowModule_1_io_V_wire_out_336 ),
       .io_V_wire_out_335( ArrayRowModule_1_io_V_wire_out_335 ),
       .io_V_wire_out_334( ArrayRowModule_1_io_V_wire_out_334 ),
       .io_V_wire_out_333( ArrayRowModule_1_io_V_wire_out_333 ),
       .io_V_wire_out_332( ArrayRowModule_1_io_V_wire_out_332 ),
       .io_V_wire_out_331( ArrayRowModule_1_io_V_wire_out_331 ),
       .io_V_wire_out_330( ArrayRowModule_1_io_V_wire_out_330 ),
       .io_V_wire_out_329( ArrayRowModule_1_io_V_wire_out_329 ),
       .io_V_wire_out_328( ArrayRowModule_1_io_V_wire_out_328 ),
       .io_V_wire_out_327( ArrayRowModule_1_io_V_wire_out_327 ),
       .io_V_wire_out_326( ArrayRowModule_1_io_V_wire_out_326 ),
       .io_V_wire_out_325( ArrayRowModule_1_io_V_wire_out_325 ),
       .io_V_wire_out_324( ArrayRowModule_1_io_V_wire_out_324 ),
       .io_V_wire_out_323( ArrayRowModule_1_io_V_wire_out_323 ),
       .io_V_wire_out_322( ArrayRowModule_1_io_V_wire_out_322 ),
       .io_V_wire_out_321( ArrayRowModule_1_io_V_wire_out_321 ),
       .io_V_wire_out_320( ArrayRowModule_1_io_V_wire_out_320 ),
       .io_V_wire_out_319( ArrayRowModule_1_io_V_wire_out_319 ),
       .io_V_wire_out_318( ArrayRowModule_1_io_V_wire_out_318 ),
       .io_V_wire_out_317( ArrayRowModule_1_io_V_wire_out_317 ),
       .io_V_wire_out_316( ArrayRowModule_1_io_V_wire_out_316 ),
       .io_V_wire_out_315( ArrayRowModule_1_io_V_wire_out_315 ),
       .io_V_wire_out_314( ArrayRowModule_1_io_V_wire_out_314 ),
       .io_V_wire_out_313( ArrayRowModule_1_io_V_wire_out_313 ),
       .io_V_wire_out_312( ArrayRowModule_1_io_V_wire_out_312 ),
       .io_V_wire_out_311( ArrayRowModule_1_io_V_wire_out_311 ),
       .io_V_wire_out_310( ArrayRowModule_1_io_V_wire_out_310 ),
       .io_V_wire_out_309( ArrayRowModule_1_io_V_wire_out_309 ),
       .io_V_wire_out_308( ArrayRowModule_1_io_V_wire_out_308 ),
       .io_V_wire_out_307( ArrayRowModule_1_io_V_wire_out_307 ),
       .io_V_wire_out_306( ArrayRowModule_1_io_V_wire_out_306 ),
       .io_V_wire_out_305( ArrayRowModule_1_io_V_wire_out_305 ),
       .io_V_wire_out_304( ArrayRowModule_1_io_V_wire_out_304 ),
       .io_V_wire_out_303( ArrayRowModule_1_io_V_wire_out_303 ),
       .io_V_wire_out_302( ArrayRowModule_1_io_V_wire_out_302 ),
       .io_V_wire_out_301( ArrayRowModule_1_io_V_wire_out_301 ),
       .io_V_wire_out_300( ArrayRowModule_1_io_V_wire_out_300 ),
       .io_V_wire_out_299( ArrayRowModule_1_io_V_wire_out_299 ),
       .io_V_wire_out_298( ArrayRowModule_1_io_V_wire_out_298 ),
       .io_V_wire_out_297( ArrayRowModule_1_io_V_wire_out_297 ),
       .io_V_wire_out_296( ArrayRowModule_1_io_V_wire_out_296 ),
       .io_V_wire_out_295( ArrayRowModule_1_io_V_wire_out_295 ),
       .io_V_wire_out_294( ArrayRowModule_1_io_V_wire_out_294 ),
       .io_V_wire_out_293( ArrayRowModule_1_io_V_wire_out_293 ),
       .io_V_wire_out_292( ArrayRowModule_1_io_V_wire_out_292 ),
       .io_V_wire_out_291( ArrayRowModule_1_io_V_wire_out_291 ),
       .io_V_wire_out_290( ArrayRowModule_1_io_V_wire_out_290 ),
       .io_V_wire_out_289( ArrayRowModule_1_io_V_wire_out_289 ),
       .io_V_wire_out_288( ArrayRowModule_1_io_V_wire_out_288 ),
       .io_V_wire_out_287( ArrayRowModule_1_io_V_wire_out_287 ),
       .io_V_wire_out_286( ArrayRowModule_1_io_V_wire_out_286 ),
       .io_V_wire_out_285( ArrayRowModule_1_io_V_wire_out_285 ),
       .io_V_wire_out_284( ArrayRowModule_1_io_V_wire_out_284 ),
       .io_V_wire_out_283( ArrayRowModule_1_io_V_wire_out_283 ),
       .io_V_wire_out_282( ArrayRowModule_1_io_V_wire_out_282 ),
       .io_V_wire_out_281( ArrayRowModule_1_io_V_wire_out_281 ),
       .io_V_wire_out_280( ArrayRowModule_1_io_V_wire_out_280 ),
       .io_V_wire_out_279( ArrayRowModule_1_io_V_wire_out_279 ),
       .io_V_wire_out_278( ArrayRowModule_1_io_V_wire_out_278 ),
       .io_V_wire_out_277( ArrayRowModule_1_io_V_wire_out_277 ),
       .io_V_wire_out_276( ArrayRowModule_1_io_V_wire_out_276 ),
       .io_V_wire_out_275( ArrayRowModule_1_io_V_wire_out_275 ),
       .io_V_wire_out_274( ArrayRowModule_1_io_V_wire_out_274 ),
       .io_V_wire_out_273( ArrayRowModule_1_io_V_wire_out_273 ),
       .io_V_wire_out_272( ArrayRowModule_1_io_V_wire_out_272 ),
       .io_V_wire_out_271( ArrayRowModule_1_io_V_wire_out_271 ),
       .io_V_wire_out_270( ArrayRowModule_1_io_V_wire_out_270 ),
       .io_V_wire_out_269( ArrayRowModule_1_io_V_wire_out_269 ),
       .io_V_wire_out_268( ArrayRowModule_1_io_V_wire_out_268 ),
       .io_V_wire_out_267( ArrayRowModule_1_io_V_wire_out_267 ),
       .io_V_wire_out_266( ArrayRowModule_1_io_V_wire_out_266 ),
       .io_V_wire_out_265( ArrayRowModule_1_io_V_wire_out_265 ),
       .io_V_wire_out_264( ArrayRowModule_1_io_V_wire_out_264 ),
       .io_V_wire_out_263( ArrayRowModule_1_io_V_wire_out_263 ),
       .io_V_wire_out_262( ArrayRowModule_1_io_V_wire_out_262 ),
       .io_V_wire_out_261( ArrayRowModule_1_io_V_wire_out_261 ),
       .io_V_wire_out_260( ArrayRowModule_1_io_V_wire_out_260 ),
       .io_V_wire_out_259( ArrayRowModule_1_io_V_wire_out_259 ),
       .io_V_wire_out_258( ArrayRowModule_1_io_V_wire_out_258 ),
       .io_V_wire_out_257( ArrayRowModule_1_io_V_wire_out_257 ),
       .io_V_wire_out_256( ArrayRowModule_1_io_V_wire_out_256 ),
       .io_V_wire_out_255( ArrayRowModule_1_io_V_wire_out_255 ),
       .io_V_wire_out_254( ArrayRowModule_1_io_V_wire_out_254 ),
       .io_V_wire_out_253( ArrayRowModule_1_io_V_wire_out_253 ),
       .io_V_wire_out_252( ArrayRowModule_1_io_V_wire_out_252 ),
       .io_V_wire_out_251( ArrayRowModule_1_io_V_wire_out_251 ),
       .io_V_wire_out_250( ArrayRowModule_1_io_V_wire_out_250 ),
       .io_V_wire_out_249( ArrayRowModule_1_io_V_wire_out_249 ),
       .io_V_wire_out_248( ArrayRowModule_1_io_V_wire_out_248 ),
       .io_V_wire_out_247( ArrayRowModule_1_io_V_wire_out_247 ),
       .io_V_wire_out_246( ArrayRowModule_1_io_V_wire_out_246 ),
       .io_V_wire_out_245( ArrayRowModule_1_io_V_wire_out_245 ),
       .io_V_wire_out_244( ArrayRowModule_1_io_V_wire_out_244 ),
       .io_V_wire_out_243( ArrayRowModule_1_io_V_wire_out_243 ),
       .io_V_wire_out_242( ArrayRowModule_1_io_V_wire_out_242 ),
       .io_V_wire_out_241( ArrayRowModule_1_io_V_wire_out_241 ),
       .io_V_wire_out_240( ArrayRowModule_1_io_V_wire_out_240 ),
       .io_V_wire_out_239( ArrayRowModule_1_io_V_wire_out_239 ),
       .io_V_wire_out_238( ArrayRowModule_1_io_V_wire_out_238 ),
       .io_V_wire_out_237( ArrayRowModule_1_io_V_wire_out_237 ),
       .io_V_wire_out_236( ArrayRowModule_1_io_V_wire_out_236 ),
       .io_V_wire_out_235( ArrayRowModule_1_io_V_wire_out_235 ),
       .io_V_wire_out_234( ArrayRowModule_1_io_V_wire_out_234 ),
       .io_V_wire_out_233( ArrayRowModule_1_io_V_wire_out_233 ),
       .io_V_wire_out_232( ArrayRowModule_1_io_V_wire_out_232 ),
       .io_V_wire_out_231( ArrayRowModule_1_io_V_wire_out_231 ),
       .io_V_wire_out_230( ArrayRowModule_1_io_V_wire_out_230 ),
       .io_V_wire_out_229( ArrayRowModule_1_io_V_wire_out_229 ),
       .io_V_wire_out_228( ArrayRowModule_1_io_V_wire_out_228 ),
       .io_V_wire_out_227( ArrayRowModule_1_io_V_wire_out_227 ),
       .io_V_wire_out_226( ArrayRowModule_1_io_V_wire_out_226 ),
       .io_V_wire_out_225( ArrayRowModule_1_io_V_wire_out_225 ),
       .io_V_wire_out_224( ArrayRowModule_1_io_V_wire_out_224 ),
       .io_V_wire_out_223( ArrayRowModule_1_io_V_wire_out_223 ),
       .io_V_wire_out_222( ArrayRowModule_1_io_V_wire_out_222 ),
       .io_V_wire_out_221( ArrayRowModule_1_io_V_wire_out_221 ),
       .io_V_wire_out_220( ArrayRowModule_1_io_V_wire_out_220 ),
       .io_V_wire_out_219( ArrayRowModule_1_io_V_wire_out_219 ),
       .io_V_wire_out_218( ArrayRowModule_1_io_V_wire_out_218 ),
       .io_V_wire_out_217( ArrayRowModule_1_io_V_wire_out_217 ),
       .io_V_wire_out_216( ArrayRowModule_1_io_V_wire_out_216 ),
       .io_V_wire_out_215( ArrayRowModule_1_io_V_wire_out_215 ),
       .io_V_wire_out_214( ArrayRowModule_1_io_V_wire_out_214 ),
       .io_V_wire_out_213( ArrayRowModule_1_io_V_wire_out_213 ),
       .io_V_wire_out_212( ArrayRowModule_1_io_V_wire_out_212 ),
       .io_V_wire_out_211( ArrayRowModule_1_io_V_wire_out_211 ),
       .io_V_wire_out_210( ArrayRowModule_1_io_V_wire_out_210 ),
       .io_V_wire_out_209( ArrayRowModule_1_io_V_wire_out_209 ),
       .io_V_wire_out_208( ArrayRowModule_1_io_V_wire_out_208 ),
       .io_V_wire_out_207( ArrayRowModule_1_io_V_wire_out_207 ),
       .io_V_wire_out_206( ArrayRowModule_1_io_V_wire_out_206 ),
       .io_V_wire_out_205( ArrayRowModule_1_io_V_wire_out_205 ),
       .io_V_wire_out_204( ArrayRowModule_1_io_V_wire_out_204 ),
       .io_V_wire_out_203( ArrayRowModule_1_io_V_wire_out_203 ),
       .io_V_wire_out_202( ArrayRowModule_1_io_V_wire_out_202 ),
       .io_V_wire_out_201( ArrayRowModule_1_io_V_wire_out_201 ),
       .io_V_wire_out_200( ArrayRowModule_1_io_V_wire_out_200 ),
       .io_V_wire_out_199( ArrayRowModule_1_io_V_wire_out_199 ),
       .io_V_wire_out_198( ArrayRowModule_1_io_V_wire_out_198 ),
       .io_V_wire_out_197( ArrayRowModule_1_io_V_wire_out_197 ),
       .io_V_wire_out_196( ArrayRowModule_1_io_V_wire_out_196 ),
       .io_V_wire_out_195( ArrayRowModule_1_io_V_wire_out_195 ),
       .io_V_wire_out_194( ArrayRowModule_1_io_V_wire_out_194 ),
       .io_V_wire_out_193( ArrayRowModule_1_io_V_wire_out_193 ),
       .io_V_wire_out_192( ArrayRowModule_1_io_V_wire_out_192 ),
       .io_V_wire_out_191( ArrayRowModule_1_io_V_wire_out_191 ),
       .io_V_wire_out_190( ArrayRowModule_1_io_V_wire_out_190 ),
       .io_V_wire_out_189( ArrayRowModule_1_io_V_wire_out_189 ),
       .io_V_wire_out_188( ArrayRowModule_1_io_V_wire_out_188 ),
       .io_V_wire_out_187( ArrayRowModule_1_io_V_wire_out_187 ),
       .io_V_wire_out_186( ArrayRowModule_1_io_V_wire_out_186 ),
       .io_V_wire_out_185( ArrayRowModule_1_io_V_wire_out_185 ),
       .io_V_wire_out_184( ArrayRowModule_1_io_V_wire_out_184 ),
       .io_V_wire_out_183( ArrayRowModule_1_io_V_wire_out_183 ),
       .io_V_wire_out_182( ArrayRowModule_1_io_V_wire_out_182 ),
       .io_V_wire_out_181( ArrayRowModule_1_io_V_wire_out_181 ),
       .io_V_wire_out_180( ArrayRowModule_1_io_V_wire_out_180 ),
       .io_V_wire_out_179( ArrayRowModule_1_io_V_wire_out_179 ),
       .io_V_wire_out_178( ArrayRowModule_1_io_V_wire_out_178 ),
       .io_V_wire_out_177( ArrayRowModule_1_io_V_wire_out_177 ),
       .io_V_wire_out_176( ArrayRowModule_1_io_V_wire_out_176 ),
       .io_V_wire_out_175( ArrayRowModule_1_io_V_wire_out_175 ),
       .io_V_wire_out_174( ArrayRowModule_1_io_V_wire_out_174 ),
       .io_V_wire_out_173( ArrayRowModule_1_io_V_wire_out_173 ),
       .io_V_wire_out_172( ArrayRowModule_1_io_V_wire_out_172 ),
       .io_V_wire_out_171( ArrayRowModule_1_io_V_wire_out_171 ),
       .io_V_wire_out_170( ArrayRowModule_1_io_V_wire_out_170 ),
       .io_V_wire_out_169( ArrayRowModule_1_io_V_wire_out_169 ),
       .io_V_wire_out_168( ArrayRowModule_1_io_V_wire_out_168 ),
       .io_V_wire_out_167( ArrayRowModule_1_io_V_wire_out_167 ),
       .io_V_wire_out_166( ArrayRowModule_1_io_V_wire_out_166 ),
       .io_V_wire_out_165( ArrayRowModule_1_io_V_wire_out_165 ),
       .io_V_wire_out_164( ArrayRowModule_1_io_V_wire_out_164 ),
       .io_V_wire_out_163( ArrayRowModule_1_io_V_wire_out_163 ),
       .io_V_wire_out_162( ArrayRowModule_1_io_V_wire_out_162 ),
       .io_V_wire_out_161( ArrayRowModule_1_io_V_wire_out_161 ),
       .io_V_wire_out_160( ArrayRowModule_1_io_V_wire_out_160 ),
       .io_V_wire_out_159( ArrayRowModule_1_io_V_wire_out_159 ),
       .io_V_wire_out_158( ArrayRowModule_1_io_V_wire_out_158 ),
       .io_V_wire_out_157( ArrayRowModule_1_io_V_wire_out_157 ),
       .io_V_wire_out_156( ArrayRowModule_1_io_V_wire_out_156 ),
       .io_V_wire_out_155( ArrayRowModule_1_io_V_wire_out_155 ),
       .io_V_wire_out_154( ArrayRowModule_1_io_V_wire_out_154 ),
       .io_V_wire_out_153( ArrayRowModule_1_io_V_wire_out_153 ),
       .io_V_wire_out_152( ArrayRowModule_1_io_V_wire_out_152 ),
       .io_V_wire_out_151( ArrayRowModule_1_io_V_wire_out_151 ),
       .io_V_wire_out_150( ArrayRowModule_1_io_V_wire_out_150 ),
       .io_V_wire_out_149( ArrayRowModule_1_io_V_wire_out_149 ),
       .io_V_wire_out_148( ArrayRowModule_1_io_V_wire_out_148 ),
       .io_V_wire_out_147( ArrayRowModule_1_io_V_wire_out_147 ),
       .io_V_wire_out_146( ArrayRowModule_1_io_V_wire_out_146 ),
       .io_V_wire_out_145( ArrayRowModule_1_io_V_wire_out_145 ),
       .io_V_wire_out_144( ArrayRowModule_1_io_V_wire_out_144 ),
       .io_V_wire_out_143( ArrayRowModule_1_io_V_wire_out_143 ),
       .io_V_wire_out_142( ArrayRowModule_1_io_V_wire_out_142 ),
       .io_V_wire_out_141( ArrayRowModule_1_io_V_wire_out_141 ),
       .io_V_wire_out_140( ArrayRowModule_1_io_V_wire_out_140 ),
       .io_V_wire_out_139( ArrayRowModule_1_io_V_wire_out_139 ),
       .io_V_wire_out_138( ArrayRowModule_1_io_V_wire_out_138 ),
       .io_V_wire_out_137( ArrayRowModule_1_io_V_wire_out_137 ),
       .io_V_wire_out_136( ArrayRowModule_1_io_V_wire_out_136 ),
       .io_V_wire_out_135( ArrayRowModule_1_io_V_wire_out_135 ),
       .io_V_wire_out_134( ArrayRowModule_1_io_V_wire_out_134 ),
       .io_V_wire_out_133( ArrayRowModule_1_io_V_wire_out_133 ),
       .io_V_wire_out_132( ArrayRowModule_1_io_V_wire_out_132 ),
       .io_V_wire_out_131( ArrayRowModule_1_io_V_wire_out_131 ),
       .io_V_wire_out_130( ArrayRowModule_1_io_V_wire_out_130 ),
       .io_V_wire_out_129( ArrayRowModule_1_io_V_wire_out_129 ),
       .io_V_wire_out_128( ArrayRowModule_1_io_V_wire_out_128 ),
       .io_V_wire_out_127( ArrayRowModule_1_io_V_wire_out_127 ),
       .io_V_wire_out_126( ArrayRowModule_1_io_V_wire_out_126 ),
       .io_V_wire_out_125( ArrayRowModule_1_io_V_wire_out_125 ),
       .io_V_wire_out_124( ArrayRowModule_1_io_V_wire_out_124 ),
       .io_V_wire_out_123( ArrayRowModule_1_io_V_wire_out_123 ),
       .io_V_wire_out_122( ArrayRowModule_1_io_V_wire_out_122 ),
       .io_V_wire_out_121( ArrayRowModule_1_io_V_wire_out_121 ),
       .io_V_wire_out_120( ArrayRowModule_1_io_V_wire_out_120 ),
       .io_V_wire_out_119( ArrayRowModule_1_io_V_wire_out_119 ),
       .io_V_wire_out_118( ArrayRowModule_1_io_V_wire_out_118 ),
       .io_V_wire_out_117( ArrayRowModule_1_io_V_wire_out_117 ),
       .io_V_wire_out_116( ArrayRowModule_1_io_V_wire_out_116 ),
       .io_V_wire_out_115( ArrayRowModule_1_io_V_wire_out_115 ),
       .io_V_wire_out_114( ArrayRowModule_1_io_V_wire_out_114 ),
       .io_V_wire_out_113( ArrayRowModule_1_io_V_wire_out_113 ),
       .io_V_wire_out_112( ArrayRowModule_1_io_V_wire_out_112 ),
       .io_V_wire_out_111( ArrayRowModule_1_io_V_wire_out_111 ),
       .io_V_wire_out_110( ArrayRowModule_1_io_V_wire_out_110 ),
       .io_V_wire_out_109( ArrayRowModule_1_io_V_wire_out_109 ),
       .io_V_wire_out_108( ArrayRowModule_1_io_V_wire_out_108 ),
       .io_V_wire_out_107( ArrayRowModule_1_io_V_wire_out_107 ),
       .io_V_wire_out_106( ArrayRowModule_1_io_V_wire_out_106 ),
       .io_V_wire_out_105( ArrayRowModule_1_io_V_wire_out_105 ),
       .io_V_wire_out_104( ArrayRowModule_1_io_V_wire_out_104 ),
       .io_V_wire_out_103( ArrayRowModule_1_io_V_wire_out_103 ),
       .io_V_wire_out_102( ArrayRowModule_1_io_V_wire_out_102 ),
       .io_V_wire_out_101( ArrayRowModule_1_io_V_wire_out_101 ),
       .io_V_wire_out_100( ArrayRowModule_1_io_V_wire_out_100 ),
       .io_V_wire_out_99( ArrayRowModule_1_io_V_wire_out_99 ),
       .io_V_wire_out_98( ArrayRowModule_1_io_V_wire_out_98 ),
       .io_V_wire_out_97( ArrayRowModule_1_io_V_wire_out_97 ),
       .io_V_wire_out_96( ArrayRowModule_1_io_V_wire_out_96 ),
       .io_V_wire_out_95( ArrayRowModule_1_io_V_wire_out_95 ),
       .io_V_wire_out_94( ArrayRowModule_1_io_V_wire_out_94 ),
       .io_V_wire_out_93( ArrayRowModule_1_io_V_wire_out_93 ),
       .io_V_wire_out_92( ArrayRowModule_1_io_V_wire_out_92 ),
       .io_V_wire_out_91( ArrayRowModule_1_io_V_wire_out_91 ),
       .io_V_wire_out_90( ArrayRowModule_1_io_V_wire_out_90 ),
       .io_V_wire_out_89( ArrayRowModule_1_io_V_wire_out_89 ),
       .io_V_wire_out_88( ArrayRowModule_1_io_V_wire_out_88 ),
       .io_V_wire_out_87( ArrayRowModule_1_io_V_wire_out_87 ),
       .io_V_wire_out_86( ArrayRowModule_1_io_V_wire_out_86 ),
       .io_V_wire_out_85( ArrayRowModule_1_io_V_wire_out_85 ),
       .io_V_wire_out_84( ArrayRowModule_1_io_V_wire_out_84 ),
       .io_V_wire_out_83( ArrayRowModule_1_io_V_wire_out_83 ),
       .io_V_wire_out_82( ArrayRowModule_1_io_V_wire_out_82 ),
       .io_V_wire_out_81( ArrayRowModule_1_io_V_wire_out_81 ),
       .io_V_wire_out_80( ArrayRowModule_1_io_V_wire_out_80 ),
       .io_V_wire_out_79( ArrayRowModule_1_io_V_wire_out_79 ),
       .io_V_wire_out_78( ArrayRowModule_1_io_V_wire_out_78 ),
       .io_V_wire_out_77( ArrayRowModule_1_io_V_wire_out_77 ),
       .io_V_wire_out_76( ArrayRowModule_1_io_V_wire_out_76 ),
       .io_V_wire_out_75( ArrayRowModule_1_io_V_wire_out_75 ),
       .io_V_wire_out_74( ArrayRowModule_1_io_V_wire_out_74 ),
       .io_V_wire_out_73( ArrayRowModule_1_io_V_wire_out_73 ),
       .io_V_wire_out_72( ArrayRowModule_1_io_V_wire_out_72 ),
       .io_V_wire_out_71( ArrayRowModule_1_io_V_wire_out_71 ),
       .io_V_wire_out_70( ArrayRowModule_1_io_V_wire_out_70 ),
       .io_V_wire_out_69( ArrayRowModule_1_io_V_wire_out_69 ),
       .io_V_wire_out_68( ArrayRowModule_1_io_V_wire_out_68 ),
       .io_V_wire_out_67( ArrayRowModule_1_io_V_wire_out_67 ),
       .io_V_wire_out_66( ArrayRowModule_1_io_V_wire_out_66 ),
       .io_V_wire_out_65( ArrayRowModule_1_io_V_wire_out_65 ),
       .io_V_wire_out_64( ArrayRowModule_1_io_V_wire_out_64 ),
       .io_V_wire_out_63( ArrayRowModule_1_io_V_wire_out_63 ),
       .io_V_wire_out_62( ArrayRowModule_1_io_V_wire_out_62 ),
       .io_V_wire_out_61( ArrayRowModule_1_io_V_wire_out_61 ),
       .io_V_wire_out_60( ArrayRowModule_1_io_V_wire_out_60 ),
       .io_V_wire_out_59( ArrayRowModule_1_io_V_wire_out_59 ),
       .io_V_wire_out_58( ArrayRowModule_1_io_V_wire_out_58 ),
       .io_V_wire_out_57( ArrayRowModule_1_io_V_wire_out_57 ),
       .io_V_wire_out_56( ArrayRowModule_1_io_V_wire_out_56 ),
       .io_V_wire_out_55( ArrayRowModule_1_io_V_wire_out_55 ),
       .io_V_wire_out_54( ArrayRowModule_1_io_V_wire_out_54 ),
       .io_V_wire_out_53( ArrayRowModule_1_io_V_wire_out_53 ),
       .io_V_wire_out_52( ArrayRowModule_1_io_V_wire_out_52 ),
       .io_V_wire_out_51( ArrayRowModule_1_io_V_wire_out_51 ),
       .io_V_wire_out_50( ArrayRowModule_1_io_V_wire_out_50 ),
       .io_V_wire_out_49( ArrayRowModule_1_io_V_wire_out_49 ),
       .io_V_wire_out_48( ArrayRowModule_1_io_V_wire_out_48 ),
       .io_V_wire_out_47( ArrayRowModule_1_io_V_wire_out_47 ),
       .io_V_wire_out_46( ArrayRowModule_1_io_V_wire_out_46 ),
       .io_V_wire_out_45( ArrayRowModule_1_io_V_wire_out_45 ),
       .io_V_wire_out_44( ArrayRowModule_1_io_V_wire_out_44 ),
       .io_V_wire_out_43( ArrayRowModule_1_io_V_wire_out_43 ),
       .io_V_wire_out_42( ArrayRowModule_1_io_V_wire_out_42 ),
       .io_V_wire_out_41( ArrayRowModule_1_io_V_wire_out_41 ),
       .io_V_wire_out_40( ArrayRowModule_1_io_V_wire_out_40 ),
       .io_V_wire_out_39( ArrayRowModule_1_io_V_wire_out_39 ),
       .io_V_wire_out_38( ArrayRowModule_1_io_V_wire_out_38 ),
       .io_V_wire_out_37( ArrayRowModule_1_io_V_wire_out_37 ),
       .io_V_wire_out_36( ArrayRowModule_1_io_V_wire_out_36 ),
       .io_V_wire_out_35( ArrayRowModule_1_io_V_wire_out_35 ),
       .io_V_wire_out_34( ArrayRowModule_1_io_V_wire_out_34 ),
       .io_V_wire_out_33( ArrayRowModule_1_io_V_wire_out_33 ),
       .io_V_wire_out_32( ArrayRowModule_1_io_V_wire_out_32 ),
       .io_V_wire_out_31( ArrayRowModule_1_io_V_wire_out_31 ),
       .io_V_wire_out_30( ArrayRowModule_1_io_V_wire_out_30 ),
       .io_V_wire_out_29( ArrayRowModule_1_io_V_wire_out_29 ),
       .io_V_wire_out_28( ArrayRowModule_1_io_V_wire_out_28 ),
       .io_V_wire_out_27( ArrayRowModule_1_io_V_wire_out_27 ),
       .io_V_wire_out_26( ArrayRowModule_1_io_V_wire_out_26 ),
       .io_V_wire_out_25( ArrayRowModule_1_io_V_wire_out_25 ),
       .io_V_wire_out_24( ArrayRowModule_1_io_V_wire_out_24 ),
       .io_V_wire_out_23( ArrayRowModule_1_io_V_wire_out_23 ),
       .io_V_wire_out_22( ArrayRowModule_1_io_V_wire_out_22 ),
       .io_V_wire_out_21( ArrayRowModule_1_io_V_wire_out_21 ),
       .io_V_wire_out_20( ArrayRowModule_1_io_V_wire_out_20 ),
       .io_V_wire_out_19( ArrayRowModule_1_io_V_wire_out_19 ),
       .io_V_wire_out_18( ArrayRowModule_1_io_V_wire_out_18 ),
       .io_V_wire_out_17( ArrayRowModule_1_io_V_wire_out_17 ),
       .io_V_wire_out_16( ArrayRowModule_1_io_V_wire_out_16 ),
       .io_V_wire_out_15( ArrayRowModule_1_io_V_wire_out_15 ),
       .io_V_wire_out_14( ArrayRowModule_1_io_V_wire_out_14 ),
       .io_V_wire_out_13( ArrayRowModule_1_io_V_wire_out_13 ),
       .io_V_wire_out_12( ArrayRowModule_1_io_V_wire_out_12 ),
       .io_V_wire_out_11( ArrayRowModule_1_io_V_wire_out_11 ),
       .io_V_wire_out_10( ArrayRowModule_1_io_V_wire_out_10 ),
       .io_V_wire_out_9( ArrayRowModule_1_io_V_wire_out_9 ),
       .io_V_wire_out_8( ArrayRowModule_1_io_V_wire_out_8 ),
       .io_V_wire_out_7( ArrayRowModule_1_io_V_wire_out_7 ),
       .io_V_wire_out_6( ArrayRowModule_1_io_V_wire_out_6 ),
       .io_V_wire_out_5( ArrayRowModule_1_io_V_wire_out_5 ),
       .io_V_wire_out_4( ArrayRowModule_1_io_V_wire_out_4 ),
       .io_V_wire_out_3( ArrayRowModule_1_io_V_wire_out_3 ),
       .io_V_wire_out_2( ArrayRowModule_1_io_V_wire_out_2 ),
       .io_V_wire_out_1( ArrayRowModule_1_io_V_wire_out_1 ),
       .io_V_wire_out_0( ArrayRowModule_1_io_V_wire_out_0 ),
       .io_V_wire_en_22( ArrayRowModule_1_io_V_wire_en_22 ),
       .io_V_wire_en_21( ArrayRowModule_1_io_V_wire_en_21 ),
       .io_V_wire_en_20( ArrayRowModule_1_io_V_wire_en_20 ),
       .io_V_wire_en_19( ArrayRowModule_1_io_V_wire_en_19 ),
       .io_V_wire_en_18( ArrayRowModule_1_io_V_wire_en_18 ),
       .io_V_wire_en_17( ArrayRowModule_1_io_V_wire_en_17 ),
       .io_V_wire_en_16( ArrayRowModule_1_io_V_wire_en_16 ),
       .io_V_wire_en_15( ArrayRowModule_1_io_V_wire_en_15 ),
       .io_V_wire_en_14( ArrayRowModule_1_io_V_wire_en_14 ),
       .io_V_wire_en_13( ArrayRowModule_1_io_V_wire_en_13 ),
       .io_V_wire_en_12( ArrayRowModule_1_io_V_wire_en_12 ),
       .io_V_wire_en_11( ArrayRowModule_1_io_V_wire_en_11 ),
       .io_V_wire_en_10( ArrayRowModule_1_io_V_wire_en_10 ),
       .io_V_wire_en_9( ArrayRowModule_1_io_V_wire_en_9 ),
       .io_V_wire_en_8( ArrayRowModule_1_io_V_wire_en_8 ),
       .io_V_wire_en_7( ArrayRowModule_1_io_V_wire_en_7 ),
       .io_V_wire_en_6( ArrayRowModule_1_io_V_wire_en_6 ),
       .io_V_wire_en_5( ArrayRowModule_1_io_V_wire_en_5 ),
       .io_V_wire_en_4( ArrayRowModule_1_io_V_wire_en_4 ),
       .io_V_wire_en_3( ArrayRowModule_1_io_V_wire_en_3 ),
       .io_V_wire_en_2( ArrayRowModule_1_io_V_wire_en_2 ),
       .io_V_wire_en_1( ArrayRowModule_1_io_V_wire_en_1 ),
       .io_V_wire_en_0( ArrayRowModule_1_io_V_wire_en_0 ),
       .io_G_wire_above_3( ArrayRowModule_io_G_wire_below_3 ),
       .io_G_wire_above_2( ArrayRowModule_io_G_wire_below_2 ),
       .io_G_wire_above_1( ArrayRowModule_io_G_wire_below_1 ),
       .io_G_wire_above_0( ArrayRowModule_io_G_wire_below_0 ),
       .io_H_wire_above_32( ArrayRowModule_io_H_wire_below_32 ),
       .io_H_wire_above_31( ArrayRowModule_io_H_wire_below_31 ),
       .io_H_wire_above_30( ArrayRowModule_io_H_wire_below_30 ),
       .io_H_wire_above_29( ArrayRowModule_io_H_wire_below_29 ),
       .io_H_wire_above_28( ArrayRowModule_io_H_wire_below_28 ),
       .io_H_wire_above_27( ArrayRowModule_io_H_wire_below_27 ),
       .io_H_wire_above_26( ArrayRowModule_io_H_wire_below_26 ),
       .io_H_wire_above_25( ArrayRowModule_io_H_wire_below_25 ),
       .io_H_wire_above_24( ArrayRowModule_io_H_wire_below_24 ),
       .io_H_wire_above_23( ArrayRowModule_io_H_wire_below_23 ),
       .io_H_wire_above_22( ArrayRowModule_io_H_wire_below_22 ),
       .io_H_wire_above_21( ArrayRowModule_io_H_wire_below_21 ),
       .io_H_wire_above_20( ArrayRowModule_io_H_wire_below_20 ),
       .io_H_wire_above_19( ArrayRowModule_io_H_wire_below_19 ),
       .io_H_wire_above_18( ArrayRowModule_io_H_wire_below_18 ),
       .io_H_wire_above_17( ArrayRowModule_io_H_wire_below_17 ),
       .io_H_wire_above_16( ArrayRowModule_io_H_wire_below_16 ),
       .io_H_wire_above_15( ArrayRowModule_io_H_wire_below_15 ),
       .io_H_wire_above_14( ArrayRowModule_io_H_wire_below_14 ),
       .io_H_wire_above_13( ArrayRowModule_io_H_wire_below_13 ),
       .io_H_wire_above_12( ArrayRowModule_io_H_wire_below_12 ),
       .io_H_wire_above_11( ArrayRowModule_io_H_wire_below_11 ),
       .io_H_wire_above_10( ArrayRowModule_io_H_wire_below_10 ),
       .io_H_wire_above_9( ArrayRowModule_io_H_wire_below_9 ),
       .io_H_wire_above_8( ArrayRowModule_io_H_wire_below_8 ),
       .io_H_wire_above_7( ArrayRowModule_io_H_wire_below_7 ),
       .io_H_wire_above_6( ArrayRowModule_io_H_wire_below_6 ),
       .io_H_wire_above_5( ArrayRowModule_io_H_wire_below_5 ),
       .io_H_wire_above_4( ArrayRowModule_io_H_wire_below_4 ),
       .io_H_wire_above_3( ArrayRowModule_io_H_wire_below_3 ),
       .io_H_wire_above_2( ArrayRowModule_io_H_wire_below_2 ),
       .io_H_wire_above_1( ArrayRowModule_io_H_wire_below_1 ),
       .io_H_wire_above_0( ArrayRowModule_io_H_wire_below_0 ),
       .io_mem_bus_in_23( ArrayRowModule_io_mem_bus_out_23 ),
       .io_mem_bus_in_22( ArrayRowModule_io_mem_bus_out_22 ),
       .io_mem_bus_in_21( ArrayRowModule_io_mem_bus_out_21 ),
       .io_mem_bus_in_20( ArrayRowModule_io_mem_bus_out_20 ),
       .io_mem_bus_in_19( ArrayRowModule_io_mem_bus_out_19 ),
       .io_mem_bus_in_18( ArrayRowModule_io_mem_bus_out_18 ),
       .io_mem_bus_in_17( ArrayRowModule_io_mem_bus_out_17 ),
       .io_mem_bus_in_16( ArrayRowModule_io_mem_bus_out_16 ),
       .io_mem_bus_in_15( ArrayRowModule_io_mem_bus_out_15 ),
       .io_mem_bus_in_14( ArrayRowModule_io_mem_bus_out_14 ),
       .io_mem_bus_in_13( ArrayRowModule_io_mem_bus_out_13 ),
       .io_mem_bus_in_12( ArrayRowModule_io_mem_bus_out_12 ),
       .io_mem_bus_in_11( ArrayRowModule_io_mem_bus_out_11 ),
       .io_mem_bus_in_10( ArrayRowModule_io_mem_bus_out_10 ),
       .io_mem_bus_in_9( ArrayRowModule_io_mem_bus_out_9 ),
       .io_mem_bus_in_8( ArrayRowModule_io_mem_bus_out_8 ),
       .io_mem_bus_in_7( ArrayRowModule_io_mem_bus_out_7 ),
       .io_mem_bus_in_6( ArrayRowModule_io_mem_bus_out_6 ),
       .io_mem_bus_in_5( ArrayRowModule_io_mem_bus_out_5 ),
       .io_mem_bus_in_4( ArrayRowModule_io_mem_bus_out_4 ),
       .io_mem_bus_in_3( ArrayRowModule_io_mem_bus_out_3 ),
       .io_mem_bus_in_2( ArrayRowModule_io_mem_bus_out_2 ),
       .io_mem_bus_in_1( ArrayRowModule_io_mem_bus_out_1 ),
       .io_mem_bus_in_0( ArrayRowModule_io_mem_bus_out_0 ),
       .io_H_out_above_22( ArrayRowModule_io_H_out_22 ),
       .io_H_out_above_21( ArrayRowModule_io_H_out_21 ),
       .io_H_out_above_20( ArrayRowModule_io_H_out_20 ),
       .io_H_out_above_19( ArrayRowModule_io_H_out_19 ),
       .io_H_out_above_18( ArrayRowModule_io_H_out_18 ),
       .io_H_out_above_17( ArrayRowModule_io_H_out_17 ),
       .io_H_out_above_16( ArrayRowModule_io_H_out_16 ),
       .io_H_out_above_15( ArrayRowModule_io_H_out_15 ),
       .io_H_out_above_14( ArrayRowModule_io_H_out_14 ),
       .io_H_out_above_13( ArrayRowModule_io_H_out_13 ),
       .io_H_out_above_12( ArrayRowModule_io_H_out_12 ),
       .io_H_out_above_11( ArrayRowModule_io_H_out_11 ),
       .io_H_out_above_10( ArrayRowModule_io_H_out_10 ),
       .io_H_out_above_9( ArrayRowModule_io_H_out_9 ),
       .io_H_out_above_8( ArrayRowModule_io_H_out_8 ),
       .io_H_out_above_7( ArrayRowModule_io_H_out_7 ),
       .io_H_out_above_6( ArrayRowModule_io_H_out_6 ),
       .io_H_out_above_5( ArrayRowModule_io_H_out_5 ),
       .io_H_out_above_4( ArrayRowModule_io_H_out_4 ),
       .io_H_out_above_3( ArrayRowModule_io_H_out_3 ),
       .io_H_out_above_2( ArrayRowModule_io_H_out_2 ),
       .io_H_out_above_1( ArrayRowModule_io_H_out_1 ),
       .io_H_out_above_0( ArrayRowModule_io_H_out_0 ),
       .io_H_out_22( ArrayRowModule_1_io_H_out_22 ),
       .io_H_out_21( ArrayRowModule_1_io_H_out_21 ),
       .io_H_out_20( ArrayRowModule_1_io_H_out_20 ),
       .io_H_out_19( ArrayRowModule_1_io_H_out_19 ),
       .io_H_out_18( ArrayRowModule_1_io_H_out_18 ),
       .io_H_out_17( ArrayRowModule_1_io_H_out_17 ),
       .io_H_out_16( ArrayRowModule_1_io_H_out_16 ),
       .io_H_out_15( ArrayRowModule_1_io_H_out_15 ),
       .io_H_out_14( ArrayRowModule_1_io_H_out_14 ),
       .io_H_out_13( ArrayRowModule_1_io_H_out_13 ),
       .io_H_out_12( ArrayRowModule_1_io_H_out_12 ),
       .io_H_out_11( ArrayRowModule_1_io_H_out_11 ),
       .io_H_out_10( ArrayRowModule_1_io_H_out_10 ),
       .io_H_out_9( ArrayRowModule_1_io_H_out_9 ),
       .io_H_out_8( ArrayRowModule_1_io_H_out_8 ),
       .io_H_out_7( ArrayRowModule_1_io_H_out_7 ),
       .io_H_out_6( ArrayRowModule_1_io_H_out_6 ),
       .io_H_out_5( ArrayRowModule_1_io_H_out_5 ),
       .io_H_out_4( ArrayRowModule_1_io_H_out_4 ),
       .io_H_out_3( ArrayRowModule_1_io_H_out_3 ),
       .io_H_out_2( ArrayRowModule_1_io_H_out_2 ),
       .io_H_out_1( ArrayRowModule_1_io_H_out_1 ),
       .io_H_out_0( ArrayRowModule_1_io_H_out_0 ),
       .io_G_wire_below_3( ArrayRowModule_1_io_G_wire_below_3 ),
       .io_G_wire_below_2( ArrayRowModule_1_io_G_wire_below_2 ),
       .io_G_wire_below_1( ArrayRowModule_1_io_G_wire_below_1 ),
       .io_G_wire_below_0( ArrayRowModule_1_io_G_wire_below_0 ),
       .io_H_wire_below_32( ArrayRowModule_1_io_H_wire_below_32 ),
       .io_H_wire_below_31( ArrayRowModule_1_io_H_wire_below_31 ),
       .io_H_wire_below_30( ArrayRowModule_1_io_H_wire_below_30 ),
       .io_H_wire_below_29( ArrayRowModule_1_io_H_wire_below_29 ),
       .io_H_wire_below_28( ArrayRowModule_1_io_H_wire_below_28 ),
       .io_H_wire_below_27( ArrayRowModule_1_io_H_wire_below_27 ),
       .io_H_wire_below_26( ArrayRowModule_1_io_H_wire_below_26 ),
       .io_H_wire_below_25( ArrayRowModule_1_io_H_wire_below_25 ),
       .io_H_wire_below_24( ArrayRowModule_1_io_H_wire_below_24 ),
       .io_H_wire_below_23( ArrayRowModule_1_io_H_wire_below_23 ),
       .io_H_wire_below_22( ArrayRowModule_1_io_H_wire_below_22 ),
       .io_H_wire_below_21( ArrayRowModule_1_io_H_wire_below_21 ),
       .io_H_wire_below_20( ArrayRowModule_1_io_H_wire_below_20 ),
       .io_H_wire_below_19( ArrayRowModule_1_io_H_wire_below_19 ),
       .io_H_wire_below_18( ArrayRowModule_1_io_H_wire_below_18 ),
       .io_H_wire_below_17( ArrayRowModule_1_io_H_wire_below_17 ),
       .io_H_wire_below_16( ArrayRowModule_1_io_H_wire_below_16 ),
       .io_H_wire_below_15( ArrayRowModule_1_io_H_wire_below_15 ),
       .io_H_wire_below_14( ArrayRowModule_1_io_H_wire_below_14 ),
       .io_H_wire_below_13( ArrayRowModule_1_io_H_wire_below_13 ),
       .io_H_wire_below_12( ArrayRowModule_1_io_H_wire_below_12 ),
       .io_H_wire_below_11( ArrayRowModule_1_io_H_wire_below_11 ),
       .io_H_wire_below_10( ArrayRowModule_1_io_H_wire_below_10 ),
       .io_H_wire_below_9( ArrayRowModule_1_io_H_wire_below_9 ),
       .io_H_wire_below_8( ArrayRowModule_1_io_H_wire_below_8 ),
       .io_H_wire_below_7( ArrayRowModule_1_io_H_wire_below_7 ),
       .io_H_wire_below_6( ArrayRowModule_1_io_H_wire_below_6 ),
       .io_H_wire_below_5( ArrayRowModule_1_io_H_wire_below_5 ),
       .io_H_wire_below_4( ArrayRowModule_1_io_H_wire_below_4 ),
       .io_H_wire_below_3( ArrayRowModule_1_io_H_wire_below_3 ),
       .io_H_wire_below_2( ArrayRowModule_1_io_H_wire_below_2 ),
       .io_H_wire_below_1( ArrayRowModule_1_io_H_wire_below_1 ),
       .io_H_wire_below_0( ArrayRowModule_1_io_H_wire_below_0 ),
       .io_row_en( T1474 ),
       //.io_config_or_load(  )
       //.io_D_or_Z(  )
       .io_mem_bus_out_23( ArrayRowModule_1_io_mem_bus_out_23 ),
       .io_mem_bus_out_22( ArrayRowModule_1_io_mem_bus_out_22 ),
       .io_mem_bus_out_21( ArrayRowModule_1_io_mem_bus_out_21 ),
       .io_mem_bus_out_20( ArrayRowModule_1_io_mem_bus_out_20 ),
       .io_mem_bus_out_19( ArrayRowModule_1_io_mem_bus_out_19 ),
       .io_mem_bus_out_18( ArrayRowModule_1_io_mem_bus_out_18 ),
       .io_mem_bus_out_17( ArrayRowModule_1_io_mem_bus_out_17 ),
       .io_mem_bus_out_16( ArrayRowModule_1_io_mem_bus_out_16 ),
       .io_mem_bus_out_15( ArrayRowModule_1_io_mem_bus_out_15 ),
       .io_mem_bus_out_14( ArrayRowModule_1_io_mem_bus_out_14 ),
       .io_mem_bus_out_13( ArrayRowModule_1_io_mem_bus_out_13 ),
       .io_mem_bus_out_12( ArrayRowModule_1_io_mem_bus_out_12 ),
       .io_mem_bus_out_11( ArrayRowModule_1_io_mem_bus_out_11 ),
       .io_mem_bus_out_10( ArrayRowModule_1_io_mem_bus_out_10 ),
       .io_mem_bus_out_9( ArrayRowModule_1_io_mem_bus_out_9 ),
       .io_mem_bus_out_8( ArrayRowModule_1_io_mem_bus_out_8 ),
       .io_mem_bus_out_7( ArrayRowModule_1_io_mem_bus_out_7 ),
       .io_mem_bus_out_6( ArrayRowModule_1_io_mem_bus_out_6 ),
       .io_mem_bus_out_5( ArrayRowModule_1_io_mem_bus_out_5 ),
       .io_mem_bus_out_4( ArrayRowModule_1_io_mem_bus_out_4 ),
       .io_mem_bus_out_3( ArrayRowModule_1_io_mem_bus_out_3 ),
       .io_mem_bus_out_2( ArrayRowModule_1_io_mem_bus_out_2 ),
       .io_mem_bus_out_1( ArrayRowModule_1_io_mem_bus_out_1 ),
       .io_mem_bus_out_0( ArrayRowModule_1_io_mem_bus_out_0 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ArrayRowModule_1.io_config_or_load = {1{$random}};
    assign ArrayRowModule_1.io_D_or_Z = {1{$random}};
    assign ArrayRowModule_1.io_mem_bus_out_23 = {1{$random}};
// synthesis translate_on
`endif
  ArrayRowModule ArrayRowModule_2(.clk(clk), .reset(reset),
       .io_V_wire_in_367( VwireModule_io_VwirePorts_2_22_15_out ),
       .io_V_wire_in_366( VwireModule_io_VwirePorts_2_22_14_out ),
       .io_V_wire_in_365( VwireModule_io_VwirePorts_2_22_13_out ),
       .io_V_wire_in_364( VwireModule_io_VwirePorts_2_22_12_out ),
       .io_V_wire_in_363( VwireModule_io_VwirePorts_2_22_11_out ),
       .io_V_wire_in_362( VwireModule_io_VwirePorts_2_22_10_out ),
       .io_V_wire_in_361( VwireModule_io_VwirePorts_2_22_9_out ),
       .io_V_wire_in_360( VwireModule_io_VwirePorts_2_22_8_out ),
       .io_V_wire_in_359( VwireModule_io_VwirePorts_2_22_7_out ),
       .io_V_wire_in_358( VwireModule_io_VwirePorts_2_22_6_out ),
       .io_V_wire_in_357( VwireModule_io_VwirePorts_2_22_5_out ),
       .io_V_wire_in_356( VwireModule_io_VwirePorts_2_22_4_out ),
       .io_V_wire_in_355( VwireModule_io_VwirePorts_2_22_3_out ),
       .io_V_wire_in_354( VwireModule_io_VwirePorts_2_22_2_out ),
       .io_V_wire_in_353( VwireModule_io_VwirePorts_2_22_1_out ),
       .io_V_wire_in_352( VwireModule_io_VwirePorts_2_22_0_out ),
       .io_V_wire_in_351( VwireModule_io_VwirePorts_2_21_15_out ),
       .io_V_wire_in_350( VwireModule_io_VwirePorts_2_21_14_out ),
       .io_V_wire_in_349( VwireModule_io_VwirePorts_2_21_13_out ),
       .io_V_wire_in_348( VwireModule_io_VwirePorts_2_21_12_out ),
       .io_V_wire_in_347( VwireModule_io_VwirePorts_2_21_11_out ),
       .io_V_wire_in_346( VwireModule_io_VwirePorts_2_21_10_out ),
       .io_V_wire_in_345( VwireModule_io_VwirePorts_2_21_9_out ),
       .io_V_wire_in_344( VwireModule_io_VwirePorts_2_21_8_out ),
       .io_V_wire_in_343( VwireModule_io_VwirePorts_2_21_7_out ),
       .io_V_wire_in_342( VwireModule_io_VwirePorts_2_21_6_out ),
       .io_V_wire_in_341( VwireModule_io_VwirePorts_2_21_5_out ),
       .io_V_wire_in_340( VwireModule_io_VwirePorts_2_21_4_out ),
       .io_V_wire_in_339( VwireModule_io_VwirePorts_2_21_3_out ),
       .io_V_wire_in_338( VwireModule_io_VwirePorts_2_21_2_out ),
       .io_V_wire_in_337( VwireModule_io_VwirePorts_2_21_1_out ),
       .io_V_wire_in_336( VwireModule_io_VwirePorts_2_21_0_out ),
       .io_V_wire_in_335( VwireModule_io_VwirePorts_2_20_15_out ),
       .io_V_wire_in_334( VwireModule_io_VwirePorts_2_20_14_out ),
       .io_V_wire_in_333( VwireModule_io_VwirePorts_2_20_13_out ),
       .io_V_wire_in_332( VwireModule_io_VwirePorts_2_20_12_out ),
       .io_V_wire_in_331( VwireModule_io_VwirePorts_2_20_11_out ),
       .io_V_wire_in_330( VwireModule_io_VwirePorts_2_20_10_out ),
       .io_V_wire_in_329( VwireModule_io_VwirePorts_2_20_9_out ),
       .io_V_wire_in_328( VwireModule_io_VwirePorts_2_20_8_out ),
       .io_V_wire_in_327( VwireModule_io_VwirePorts_2_20_7_out ),
       .io_V_wire_in_326( VwireModule_io_VwirePorts_2_20_6_out ),
       .io_V_wire_in_325( VwireModule_io_VwirePorts_2_20_5_out ),
       .io_V_wire_in_324( VwireModule_io_VwirePorts_2_20_4_out ),
       .io_V_wire_in_323( VwireModule_io_VwirePorts_2_20_3_out ),
       .io_V_wire_in_322( VwireModule_io_VwirePorts_2_20_2_out ),
       .io_V_wire_in_321( VwireModule_io_VwirePorts_2_20_1_out ),
       .io_V_wire_in_320( VwireModule_io_VwirePorts_2_20_0_out ),
       .io_V_wire_in_319( VwireModule_io_VwirePorts_2_19_15_out ),
       .io_V_wire_in_318( VwireModule_io_VwirePorts_2_19_14_out ),
       .io_V_wire_in_317( VwireModule_io_VwirePorts_2_19_13_out ),
       .io_V_wire_in_316( VwireModule_io_VwirePorts_2_19_12_out ),
       .io_V_wire_in_315( VwireModule_io_VwirePorts_2_19_11_out ),
       .io_V_wire_in_314( VwireModule_io_VwirePorts_2_19_10_out ),
       .io_V_wire_in_313( VwireModule_io_VwirePorts_2_19_9_out ),
       .io_V_wire_in_312( VwireModule_io_VwirePorts_2_19_8_out ),
       .io_V_wire_in_311( VwireModule_io_VwirePorts_2_19_7_out ),
       .io_V_wire_in_310( VwireModule_io_VwirePorts_2_19_6_out ),
       .io_V_wire_in_309( VwireModule_io_VwirePorts_2_19_5_out ),
       .io_V_wire_in_308( VwireModule_io_VwirePorts_2_19_4_out ),
       .io_V_wire_in_307( VwireModule_io_VwirePorts_2_19_3_out ),
       .io_V_wire_in_306( VwireModule_io_VwirePorts_2_19_2_out ),
       .io_V_wire_in_305( VwireModule_io_VwirePorts_2_19_1_out ),
       .io_V_wire_in_304( VwireModule_io_VwirePorts_2_19_0_out ),
       .io_V_wire_in_303( VwireModule_io_VwirePorts_2_18_15_out ),
       .io_V_wire_in_302( VwireModule_io_VwirePorts_2_18_14_out ),
       .io_V_wire_in_301( VwireModule_io_VwirePorts_2_18_13_out ),
       .io_V_wire_in_300( VwireModule_io_VwirePorts_2_18_12_out ),
       .io_V_wire_in_299( VwireModule_io_VwirePorts_2_18_11_out ),
       .io_V_wire_in_298( VwireModule_io_VwirePorts_2_18_10_out ),
       .io_V_wire_in_297( VwireModule_io_VwirePorts_2_18_9_out ),
       .io_V_wire_in_296( VwireModule_io_VwirePorts_2_18_8_out ),
       .io_V_wire_in_295( VwireModule_io_VwirePorts_2_18_7_out ),
       .io_V_wire_in_294( VwireModule_io_VwirePorts_2_18_6_out ),
       .io_V_wire_in_293( VwireModule_io_VwirePorts_2_18_5_out ),
       .io_V_wire_in_292( VwireModule_io_VwirePorts_2_18_4_out ),
       .io_V_wire_in_291( VwireModule_io_VwirePorts_2_18_3_out ),
       .io_V_wire_in_290( VwireModule_io_VwirePorts_2_18_2_out ),
       .io_V_wire_in_289( VwireModule_io_VwirePorts_2_18_1_out ),
       .io_V_wire_in_288( VwireModule_io_VwirePorts_2_18_0_out ),
       .io_V_wire_in_287( VwireModule_io_VwirePorts_2_17_15_out ),
       .io_V_wire_in_286( VwireModule_io_VwirePorts_2_17_14_out ),
       .io_V_wire_in_285( VwireModule_io_VwirePorts_2_17_13_out ),
       .io_V_wire_in_284( VwireModule_io_VwirePorts_2_17_12_out ),
       .io_V_wire_in_283( VwireModule_io_VwirePorts_2_17_11_out ),
       .io_V_wire_in_282( VwireModule_io_VwirePorts_2_17_10_out ),
       .io_V_wire_in_281( VwireModule_io_VwirePorts_2_17_9_out ),
       .io_V_wire_in_280( VwireModule_io_VwirePorts_2_17_8_out ),
       .io_V_wire_in_279( VwireModule_io_VwirePorts_2_17_7_out ),
       .io_V_wire_in_278( VwireModule_io_VwirePorts_2_17_6_out ),
       .io_V_wire_in_277( VwireModule_io_VwirePorts_2_17_5_out ),
       .io_V_wire_in_276( VwireModule_io_VwirePorts_2_17_4_out ),
       .io_V_wire_in_275( VwireModule_io_VwirePorts_2_17_3_out ),
       .io_V_wire_in_274( VwireModule_io_VwirePorts_2_17_2_out ),
       .io_V_wire_in_273( VwireModule_io_VwirePorts_2_17_1_out ),
       .io_V_wire_in_272( VwireModule_io_VwirePorts_2_17_0_out ),
       .io_V_wire_in_271( VwireModule_io_VwirePorts_2_16_15_out ),
       .io_V_wire_in_270( VwireModule_io_VwirePorts_2_16_14_out ),
       .io_V_wire_in_269( VwireModule_io_VwirePorts_2_16_13_out ),
       .io_V_wire_in_268( VwireModule_io_VwirePorts_2_16_12_out ),
       .io_V_wire_in_267( VwireModule_io_VwirePorts_2_16_11_out ),
       .io_V_wire_in_266( VwireModule_io_VwirePorts_2_16_10_out ),
       .io_V_wire_in_265( VwireModule_io_VwirePorts_2_16_9_out ),
       .io_V_wire_in_264( VwireModule_io_VwirePorts_2_16_8_out ),
       .io_V_wire_in_263( VwireModule_io_VwirePorts_2_16_7_out ),
       .io_V_wire_in_262( VwireModule_io_VwirePorts_2_16_6_out ),
       .io_V_wire_in_261( VwireModule_io_VwirePorts_2_16_5_out ),
       .io_V_wire_in_260( VwireModule_io_VwirePorts_2_16_4_out ),
       .io_V_wire_in_259( VwireModule_io_VwirePorts_2_16_3_out ),
       .io_V_wire_in_258( VwireModule_io_VwirePorts_2_16_2_out ),
       .io_V_wire_in_257( VwireModule_io_VwirePorts_2_16_1_out ),
       .io_V_wire_in_256( VwireModule_io_VwirePorts_2_16_0_out ),
       .io_V_wire_in_255( VwireModule_io_VwirePorts_2_15_15_out ),
       .io_V_wire_in_254( VwireModule_io_VwirePorts_2_15_14_out ),
       .io_V_wire_in_253( VwireModule_io_VwirePorts_2_15_13_out ),
       .io_V_wire_in_252( VwireModule_io_VwirePorts_2_15_12_out ),
       .io_V_wire_in_251( VwireModule_io_VwirePorts_2_15_11_out ),
       .io_V_wire_in_250( VwireModule_io_VwirePorts_2_15_10_out ),
       .io_V_wire_in_249( VwireModule_io_VwirePorts_2_15_9_out ),
       .io_V_wire_in_248( VwireModule_io_VwirePorts_2_15_8_out ),
       .io_V_wire_in_247( VwireModule_io_VwirePorts_2_15_7_out ),
       .io_V_wire_in_246( VwireModule_io_VwirePorts_2_15_6_out ),
       .io_V_wire_in_245( VwireModule_io_VwirePorts_2_15_5_out ),
       .io_V_wire_in_244( VwireModule_io_VwirePorts_2_15_4_out ),
       .io_V_wire_in_243( VwireModule_io_VwirePorts_2_15_3_out ),
       .io_V_wire_in_242( VwireModule_io_VwirePorts_2_15_2_out ),
       .io_V_wire_in_241( VwireModule_io_VwirePorts_2_15_1_out ),
       .io_V_wire_in_240( VwireModule_io_VwirePorts_2_15_0_out ),
       .io_V_wire_in_239( VwireModule_io_VwirePorts_2_14_15_out ),
       .io_V_wire_in_238( VwireModule_io_VwirePorts_2_14_14_out ),
       .io_V_wire_in_237( VwireModule_io_VwirePorts_2_14_13_out ),
       .io_V_wire_in_236( VwireModule_io_VwirePorts_2_14_12_out ),
       .io_V_wire_in_235( VwireModule_io_VwirePorts_2_14_11_out ),
       .io_V_wire_in_234( VwireModule_io_VwirePorts_2_14_10_out ),
       .io_V_wire_in_233( VwireModule_io_VwirePorts_2_14_9_out ),
       .io_V_wire_in_232( VwireModule_io_VwirePorts_2_14_8_out ),
       .io_V_wire_in_231( VwireModule_io_VwirePorts_2_14_7_out ),
       .io_V_wire_in_230( VwireModule_io_VwirePorts_2_14_6_out ),
       .io_V_wire_in_229( VwireModule_io_VwirePorts_2_14_5_out ),
       .io_V_wire_in_228( VwireModule_io_VwirePorts_2_14_4_out ),
       .io_V_wire_in_227( VwireModule_io_VwirePorts_2_14_3_out ),
       .io_V_wire_in_226( VwireModule_io_VwirePorts_2_14_2_out ),
       .io_V_wire_in_225( VwireModule_io_VwirePorts_2_14_1_out ),
       .io_V_wire_in_224( VwireModule_io_VwirePorts_2_14_0_out ),
       .io_V_wire_in_223( VwireModule_io_VwirePorts_2_13_15_out ),
       .io_V_wire_in_222( VwireModule_io_VwirePorts_2_13_14_out ),
       .io_V_wire_in_221( VwireModule_io_VwirePorts_2_13_13_out ),
       .io_V_wire_in_220( VwireModule_io_VwirePorts_2_13_12_out ),
       .io_V_wire_in_219( VwireModule_io_VwirePorts_2_13_11_out ),
       .io_V_wire_in_218( VwireModule_io_VwirePorts_2_13_10_out ),
       .io_V_wire_in_217( VwireModule_io_VwirePorts_2_13_9_out ),
       .io_V_wire_in_216( VwireModule_io_VwirePorts_2_13_8_out ),
       .io_V_wire_in_215( VwireModule_io_VwirePorts_2_13_7_out ),
       .io_V_wire_in_214( VwireModule_io_VwirePorts_2_13_6_out ),
       .io_V_wire_in_213( VwireModule_io_VwirePorts_2_13_5_out ),
       .io_V_wire_in_212( VwireModule_io_VwirePorts_2_13_4_out ),
       .io_V_wire_in_211( VwireModule_io_VwirePorts_2_13_3_out ),
       .io_V_wire_in_210( VwireModule_io_VwirePorts_2_13_2_out ),
       .io_V_wire_in_209( VwireModule_io_VwirePorts_2_13_1_out ),
       .io_V_wire_in_208( VwireModule_io_VwirePorts_2_13_0_out ),
       .io_V_wire_in_207( VwireModule_io_VwirePorts_2_12_15_out ),
       .io_V_wire_in_206( VwireModule_io_VwirePorts_2_12_14_out ),
       .io_V_wire_in_205( VwireModule_io_VwirePorts_2_12_13_out ),
       .io_V_wire_in_204( VwireModule_io_VwirePorts_2_12_12_out ),
       .io_V_wire_in_203( VwireModule_io_VwirePorts_2_12_11_out ),
       .io_V_wire_in_202( VwireModule_io_VwirePorts_2_12_10_out ),
       .io_V_wire_in_201( VwireModule_io_VwirePorts_2_12_9_out ),
       .io_V_wire_in_200( VwireModule_io_VwirePorts_2_12_8_out ),
       .io_V_wire_in_199( VwireModule_io_VwirePorts_2_12_7_out ),
       .io_V_wire_in_198( VwireModule_io_VwirePorts_2_12_6_out ),
       .io_V_wire_in_197( VwireModule_io_VwirePorts_2_12_5_out ),
       .io_V_wire_in_196( VwireModule_io_VwirePorts_2_12_4_out ),
       .io_V_wire_in_195( VwireModule_io_VwirePorts_2_12_3_out ),
       .io_V_wire_in_194( VwireModule_io_VwirePorts_2_12_2_out ),
       .io_V_wire_in_193( VwireModule_io_VwirePorts_2_12_1_out ),
       .io_V_wire_in_192( VwireModule_io_VwirePorts_2_12_0_out ),
       .io_V_wire_in_191( VwireModule_io_VwirePorts_2_11_15_out ),
       .io_V_wire_in_190( VwireModule_io_VwirePorts_2_11_14_out ),
       .io_V_wire_in_189( VwireModule_io_VwirePorts_2_11_13_out ),
       .io_V_wire_in_188( VwireModule_io_VwirePorts_2_11_12_out ),
       .io_V_wire_in_187( VwireModule_io_VwirePorts_2_11_11_out ),
       .io_V_wire_in_186( VwireModule_io_VwirePorts_2_11_10_out ),
       .io_V_wire_in_185( VwireModule_io_VwirePorts_2_11_9_out ),
       .io_V_wire_in_184( VwireModule_io_VwirePorts_2_11_8_out ),
       .io_V_wire_in_183( VwireModule_io_VwirePorts_2_11_7_out ),
       .io_V_wire_in_182( VwireModule_io_VwirePorts_2_11_6_out ),
       .io_V_wire_in_181( VwireModule_io_VwirePorts_2_11_5_out ),
       .io_V_wire_in_180( VwireModule_io_VwirePorts_2_11_4_out ),
       .io_V_wire_in_179( VwireModule_io_VwirePorts_2_11_3_out ),
       .io_V_wire_in_178( VwireModule_io_VwirePorts_2_11_2_out ),
       .io_V_wire_in_177( VwireModule_io_VwirePorts_2_11_1_out ),
       .io_V_wire_in_176( VwireModule_io_VwirePorts_2_11_0_out ),
       .io_V_wire_in_175( VwireModule_io_VwirePorts_2_10_15_out ),
       .io_V_wire_in_174( VwireModule_io_VwirePorts_2_10_14_out ),
       .io_V_wire_in_173( VwireModule_io_VwirePorts_2_10_13_out ),
       .io_V_wire_in_172( VwireModule_io_VwirePorts_2_10_12_out ),
       .io_V_wire_in_171( VwireModule_io_VwirePorts_2_10_11_out ),
       .io_V_wire_in_170( VwireModule_io_VwirePorts_2_10_10_out ),
       .io_V_wire_in_169( VwireModule_io_VwirePorts_2_10_9_out ),
       .io_V_wire_in_168( VwireModule_io_VwirePorts_2_10_8_out ),
       .io_V_wire_in_167( VwireModule_io_VwirePorts_2_10_7_out ),
       .io_V_wire_in_166( VwireModule_io_VwirePorts_2_10_6_out ),
       .io_V_wire_in_165( VwireModule_io_VwirePorts_2_10_5_out ),
       .io_V_wire_in_164( VwireModule_io_VwirePorts_2_10_4_out ),
       .io_V_wire_in_163( VwireModule_io_VwirePorts_2_10_3_out ),
       .io_V_wire_in_162( VwireModule_io_VwirePorts_2_10_2_out ),
       .io_V_wire_in_161( VwireModule_io_VwirePorts_2_10_1_out ),
       .io_V_wire_in_160( VwireModule_io_VwirePorts_2_10_0_out ),
       .io_V_wire_in_159( VwireModule_io_VwirePorts_2_9_15_out ),
       .io_V_wire_in_158( VwireModule_io_VwirePorts_2_9_14_out ),
       .io_V_wire_in_157( VwireModule_io_VwirePorts_2_9_13_out ),
       .io_V_wire_in_156( VwireModule_io_VwirePorts_2_9_12_out ),
       .io_V_wire_in_155( VwireModule_io_VwirePorts_2_9_11_out ),
       .io_V_wire_in_154( VwireModule_io_VwirePorts_2_9_10_out ),
       .io_V_wire_in_153( VwireModule_io_VwirePorts_2_9_9_out ),
       .io_V_wire_in_152( VwireModule_io_VwirePorts_2_9_8_out ),
       .io_V_wire_in_151( VwireModule_io_VwirePorts_2_9_7_out ),
       .io_V_wire_in_150( VwireModule_io_VwirePorts_2_9_6_out ),
       .io_V_wire_in_149( VwireModule_io_VwirePorts_2_9_5_out ),
       .io_V_wire_in_148( VwireModule_io_VwirePorts_2_9_4_out ),
       .io_V_wire_in_147( VwireModule_io_VwirePorts_2_9_3_out ),
       .io_V_wire_in_146( VwireModule_io_VwirePorts_2_9_2_out ),
       .io_V_wire_in_145( VwireModule_io_VwirePorts_2_9_1_out ),
       .io_V_wire_in_144( VwireModule_io_VwirePorts_2_9_0_out ),
       .io_V_wire_in_143( VwireModule_io_VwirePorts_2_8_15_out ),
       .io_V_wire_in_142( VwireModule_io_VwirePorts_2_8_14_out ),
       .io_V_wire_in_141( VwireModule_io_VwirePorts_2_8_13_out ),
       .io_V_wire_in_140( VwireModule_io_VwirePorts_2_8_12_out ),
       .io_V_wire_in_139( VwireModule_io_VwirePorts_2_8_11_out ),
       .io_V_wire_in_138( VwireModule_io_VwirePorts_2_8_10_out ),
       .io_V_wire_in_137( VwireModule_io_VwirePorts_2_8_9_out ),
       .io_V_wire_in_136( VwireModule_io_VwirePorts_2_8_8_out ),
       .io_V_wire_in_135( VwireModule_io_VwirePorts_2_8_7_out ),
       .io_V_wire_in_134( VwireModule_io_VwirePorts_2_8_6_out ),
       .io_V_wire_in_133( VwireModule_io_VwirePorts_2_8_5_out ),
       .io_V_wire_in_132( VwireModule_io_VwirePorts_2_8_4_out ),
       .io_V_wire_in_131( VwireModule_io_VwirePorts_2_8_3_out ),
       .io_V_wire_in_130( VwireModule_io_VwirePorts_2_8_2_out ),
       .io_V_wire_in_129( VwireModule_io_VwirePorts_2_8_1_out ),
       .io_V_wire_in_128( VwireModule_io_VwirePorts_2_8_0_out ),
       .io_V_wire_in_127( VwireModule_io_VwirePorts_2_7_15_out ),
       .io_V_wire_in_126( VwireModule_io_VwirePorts_2_7_14_out ),
       .io_V_wire_in_125( VwireModule_io_VwirePorts_2_7_13_out ),
       .io_V_wire_in_124( VwireModule_io_VwirePorts_2_7_12_out ),
       .io_V_wire_in_123( VwireModule_io_VwirePorts_2_7_11_out ),
       .io_V_wire_in_122( VwireModule_io_VwirePorts_2_7_10_out ),
       .io_V_wire_in_121( VwireModule_io_VwirePorts_2_7_9_out ),
       .io_V_wire_in_120( VwireModule_io_VwirePorts_2_7_8_out ),
       .io_V_wire_in_119( VwireModule_io_VwirePorts_2_7_7_out ),
       .io_V_wire_in_118( VwireModule_io_VwirePorts_2_7_6_out ),
       .io_V_wire_in_117( VwireModule_io_VwirePorts_2_7_5_out ),
       .io_V_wire_in_116( VwireModule_io_VwirePorts_2_7_4_out ),
       .io_V_wire_in_115( VwireModule_io_VwirePorts_2_7_3_out ),
       .io_V_wire_in_114( VwireModule_io_VwirePorts_2_7_2_out ),
       .io_V_wire_in_113( VwireModule_io_VwirePorts_2_7_1_out ),
       .io_V_wire_in_112( VwireModule_io_VwirePorts_2_7_0_out ),
       .io_V_wire_in_111( VwireModule_io_VwirePorts_2_6_15_out ),
       .io_V_wire_in_110( VwireModule_io_VwirePorts_2_6_14_out ),
       .io_V_wire_in_109( VwireModule_io_VwirePorts_2_6_13_out ),
       .io_V_wire_in_108( VwireModule_io_VwirePorts_2_6_12_out ),
       .io_V_wire_in_107( VwireModule_io_VwirePorts_2_6_11_out ),
       .io_V_wire_in_106( VwireModule_io_VwirePorts_2_6_10_out ),
       .io_V_wire_in_105( VwireModule_io_VwirePorts_2_6_9_out ),
       .io_V_wire_in_104( VwireModule_io_VwirePorts_2_6_8_out ),
       .io_V_wire_in_103( VwireModule_io_VwirePorts_2_6_7_out ),
       .io_V_wire_in_102( VwireModule_io_VwirePorts_2_6_6_out ),
       .io_V_wire_in_101( VwireModule_io_VwirePorts_2_6_5_out ),
       .io_V_wire_in_100( VwireModule_io_VwirePorts_2_6_4_out ),
       .io_V_wire_in_99( VwireModule_io_VwirePorts_2_6_3_out ),
       .io_V_wire_in_98( VwireModule_io_VwirePorts_2_6_2_out ),
       .io_V_wire_in_97( VwireModule_io_VwirePorts_2_6_1_out ),
       .io_V_wire_in_96( VwireModule_io_VwirePorts_2_6_0_out ),
       .io_V_wire_in_95( VwireModule_io_VwirePorts_2_5_15_out ),
       .io_V_wire_in_94( VwireModule_io_VwirePorts_2_5_14_out ),
       .io_V_wire_in_93( VwireModule_io_VwirePorts_2_5_13_out ),
       .io_V_wire_in_92( VwireModule_io_VwirePorts_2_5_12_out ),
       .io_V_wire_in_91( VwireModule_io_VwirePorts_2_5_11_out ),
       .io_V_wire_in_90( VwireModule_io_VwirePorts_2_5_10_out ),
       .io_V_wire_in_89( VwireModule_io_VwirePorts_2_5_9_out ),
       .io_V_wire_in_88( VwireModule_io_VwirePorts_2_5_8_out ),
       .io_V_wire_in_87( VwireModule_io_VwirePorts_2_5_7_out ),
       .io_V_wire_in_86( VwireModule_io_VwirePorts_2_5_6_out ),
       .io_V_wire_in_85( VwireModule_io_VwirePorts_2_5_5_out ),
       .io_V_wire_in_84( VwireModule_io_VwirePorts_2_5_4_out ),
       .io_V_wire_in_83( VwireModule_io_VwirePorts_2_5_3_out ),
       .io_V_wire_in_82( VwireModule_io_VwirePorts_2_5_2_out ),
       .io_V_wire_in_81( VwireModule_io_VwirePorts_2_5_1_out ),
       .io_V_wire_in_80( VwireModule_io_VwirePorts_2_5_0_out ),
       .io_V_wire_in_79( VwireModule_io_VwirePorts_2_4_15_out ),
       .io_V_wire_in_78( VwireModule_io_VwirePorts_2_4_14_out ),
       .io_V_wire_in_77( VwireModule_io_VwirePorts_2_4_13_out ),
       .io_V_wire_in_76( VwireModule_io_VwirePorts_2_4_12_out ),
       .io_V_wire_in_75( VwireModule_io_VwirePorts_2_4_11_out ),
       .io_V_wire_in_74( VwireModule_io_VwirePorts_2_4_10_out ),
       .io_V_wire_in_73( VwireModule_io_VwirePorts_2_4_9_out ),
       .io_V_wire_in_72( VwireModule_io_VwirePorts_2_4_8_out ),
       .io_V_wire_in_71( VwireModule_io_VwirePorts_2_4_7_out ),
       .io_V_wire_in_70( VwireModule_io_VwirePorts_2_4_6_out ),
       .io_V_wire_in_69( VwireModule_io_VwirePorts_2_4_5_out ),
       .io_V_wire_in_68( VwireModule_io_VwirePorts_2_4_4_out ),
       .io_V_wire_in_67( VwireModule_io_VwirePorts_2_4_3_out ),
       .io_V_wire_in_66( VwireModule_io_VwirePorts_2_4_2_out ),
       .io_V_wire_in_65( VwireModule_io_VwirePorts_2_4_1_out ),
       .io_V_wire_in_64( VwireModule_io_VwirePorts_2_4_0_out ),
       .io_V_wire_in_63( VwireModule_io_VwirePorts_2_3_15_out ),
       .io_V_wire_in_62( VwireModule_io_VwirePorts_2_3_14_out ),
       .io_V_wire_in_61( VwireModule_io_VwirePorts_2_3_13_out ),
       .io_V_wire_in_60( VwireModule_io_VwirePorts_2_3_12_out ),
       .io_V_wire_in_59( VwireModule_io_VwirePorts_2_3_11_out ),
       .io_V_wire_in_58( VwireModule_io_VwirePorts_2_3_10_out ),
       .io_V_wire_in_57( VwireModule_io_VwirePorts_2_3_9_out ),
       .io_V_wire_in_56( VwireModule_io_VwirePorts_2_3_8_out ),
       .io_V_wire_in_55( VwireModule_io_VwirePorts_2_3_7_out ),
       .io_V_wire_in_54( VwireModule_io_VwirePorts_2_3_6_out ),
       .io_V_wire_in_53( VwireModule_io_VwirePorts_2_3_5_out ),
       .io_V_wire_in_52( VwireModule_io_VwirePorts_2_3_4_out ),
       .io_V_wire_in_51( VwireModule_io_VwirePorts_2_3_3_out ),
       .io_V_wire_in_50( VwireModule_io_VwirePorts_2_3_2_out ),
       .io_V_wire_in_49( VwireModule_io_VwirePorts_2_3_1_out ),
       .io_V_wire_in_48( VwireModule_io_VwirePorts_2_3_0_out ),
       .io_V_wire_in_47( VwireModule_io_VwirePorts_2_2_15_out ),
       .io_V_wire_in_46( VwireModule_io_VwirePorts_2_2_14_out ),
       .io_V_wire_in_45( VwireModule_io_VwirePorts_2_2_13_out ),
       .io_V_wire_in_44( VwireModule_io_VwirePorts_2_2_12_out ),
       .io_V_wire_in_43( VwireModule_io_VwirePorts_2_2_11_out ),
       .io_V_wire_in_42( VwireModule_io_VwirePorts_2_2_10_out ),
       .io_V_wire_in_41( VwireModule_io_VwirePorts_2_2_9_out ),
       .io_V_wire_in_40( VwireModule_io_VwirePorts_2_2_8_out ),
       .io_V_wire_in_39( VwireModule_io_VwirePorts_2_2_7_out ),
       .io_V_wire_in_38( VwireModule_io_VwirePorts_2_2_6_out ),
       .io_V_wire_in_37( VwireModule_io_VwirePorts_2_2_5_out ),
       .io_V_wire_in_36( VwireModule_io_VwirePorts_2_2_4_out ),
       .io_V_wire_in_35( VwireModule_io_VwirePorts_2_2_3_out ),
       .io_V_wire_in_34( VwireModule_io_VwirePorts_2_2_2_out ),
       .io_V_wire_in_33( VwireModule_io_VwirePorts_2_2_1_out ),
       .io_V_wire_in_32( VwireModule_io_VwirePorts_2_2_0_out ),
       .io_V_wire_in_31( VwireModule_io_VwirePorts_2_1_15_out ),
       .io_V_wire_in_30( VwireModule_io_VwirePorts_2_1_14_out ),
       .io_V_wire_in_29( VwireModule_io_VwirePorts_2_1_13_out ),
       .io_V_wire_in_28( VwireModule_io_VwirePorts_2_1_12_out ),
       .io_V_wire_in_27( VwireModule_io_VwirePorts_2_1_11_out ),
       .io_V_wire_in_26( VwireModule_io_VwirePorts_2_1_10_out ),
       .io_V_wire_in_25( VwireModule_io_VwirePorts_2_1_9_out ),
       .io_V_wire_in_24( VwireModule_io_VwirePorts_2_1_8_out ),
       .io_V_wire_in_23( VwireModule_io_VwirePorts_2_1_7_out ),
       .io_V_wire_in_22( VwireModule_io_VwirePorts_2_1_6_out ),
       .io_V_wire_in_21( VwireModule_io_VwirePorts_2_1_5_out ),
       .io_V_wire_in_20( VwireModule_io_VwirePorts_2_1_4_out ),
       .io_V_wire_in_19( VwireModule_io_VwirePorts_2_1_3_out ),
       .io_V_wire_in_18( VwireModule_io_VwirePorts_2_1_2_out ),
       .io_V_wire_in_17( VwireModule_io_VwirePorts_2_1_1_out ),
       .io_V_wire_in_16( VwireModule_io_VwirePorts_2_1_0_out ),
       .io_V_wire_in_15( VwireModule_io_VwirePorts_2_0_15_out ),
       .io_V_wire_in_14( VwireModule_io_VwirePorts_2_0_14_out ),
       .io_V_wire_in_13( VwireModule_io_VwirePorts_2_0_13_out ),
       .io_V_wire_in_12( VwireModule_io_VwirePorts_2_0_12_out ),
       .io_V_wire_in_11( VwireModule_io_VwirePorts_2_0_11_out ),
       .io_V_wire_in_10( VwireModule_io_VwirePorts_2_0_10_out ),
       .io_V_wire_in_9( VwireModule_io_VwirePorts_2_0_9_out ),
       .io_V_wire_in_8( VwireModule_io_VwirePorts_2_0_8_out ),
       .io_V_wire_in_7( VwireModule_io_VwirePorts_2_0_7_out ),
       .io_V_wire_in_6( VwireModule_io_VwirePorts_2_0_6_out ),
       .io_V_wire_in_5( VwireModule_io_VwirePorts_2_0_5_out ),
       .io_V_wire_in_4( VwireModule_io_VwirePorts_2_0_4_out ),
       .io_V_wire_in_3( VwireModule_io_VwirePorts_2_0_3_out ),
       .io_V_wire_in_2( VwireModule_io_VwirePorts_2_0_2_out ),
       .io_V_wire_in_1( VwireModule_io_VwirePorts_2_0_1_out ),
       .io_V_wire_in_0( VwireModule_io_VwirePorts_2_0_0_out ),
       .io_V_wire_out_367( ArrayRowModule_2_io_V_wire_out_367 ),
       .io_V_wire_out_366( ArrayRowModule_2_io_V_wire_out_366 ),
       .io_V_wire_out_365( ArrayRowModule_2_io_V_wire_out_365 ),
       .io_V_wire_out_364( ArrayRowModule_2_io_V_wire_out_364 ),
       .io_V_wire_out_363( ArrayRowModule_2_io_V_wire_out_363 ),
       .io_V_wire_out_362( ArrayRowModule_2_io_V_wire_out_362 ),
       .io_V_wire_out_361( ArrayRowModule_2_io_V_wire_out_361 ),
       .io_V_wire_out_360( ArrayRowModule_2_io_V_wire_out_360 ),
       .io_V_wire_out_359( ArrayRowModule_2_io_V_wire_out_359 ),
       .io_V_wire_out_358( ArrayRowModule_2_io_V_wire_out_358 ),
       .io_V_wire_out_357( ArrayRowModule_2_io_V_wire_out_357 ),
       .io_V_wire_out_356( ArrayRowModule_2_io_V_wire_out_356 ),
       .io_V_wire_out_355( ArrayRowModule_2_io_V_wire_out_355 ),
       .io_V_wire_out_354( ArrayRowModule_2_io_V_wire_out_354 ),
       .io_V_wire_out_353( ArrayRowModule_2_io_V_wire_out_353 ),
       .io_V_wire_out_352( ArrayRowModule_2_io_V_wire_out_352 ),
       .io_V_wire_out_351( ArrayRowModule_2_io_V_wire_out_351 ),
       .io_V_wire_out_350( ArrayRowModule_2_io_V_wire_out_350 ),
       .io_V_wire_out_349( ArrayRowModule_2_io_V_wire_out_349 ),
       .io_V_wire_out_348( ArrayRowModule_2_io_V_wire_out_348 ),
       .io_V_wire_out_347( ArrayRowModule_2_io_V_wire_out_347 ),
       .io_V_wire_out_346( ArrayRowModule_2_io_V_wire_out_346 ),
       .io_V_wire_out_345( ArrayRowModule_2_io_V_wire_out_345 ),
       .io_V_wire_out_344( ArrayRowModule_2_io_V_wire_out_344 ),
       .io_V_wire_out_343( ArrayRowModule_2_io_V_wire_out_343 ),
       .io_V_wire_out_342( ArrayRowModule_2_io_V_wire_out_342 ),
       .io_V_wire_out_341( ArrayRowModule_2_io_V_wire_out_341 ),
       .io_V_wire_out_340( ArrayRowModule_2_io_V_wire_out_340 ),
       .io_V_wire_out_339( ArrayRowModule_2_io_V_wire_out_339 ),
       .io_V_wire_out_338( ArrayRowModule_2_io_V_wire_out_338 ),
       .io_V_wire_out_337( ArrayRowModule_2_io_V_wire_out_337 ),
       .io_V_wire_out_336( ArrayRowModule_2_io_V_wire_out_336 ),
       .io_V_wire_out_335( ArrayRowModule_2_io_V_wire_out_335 ),
       .io_V_wire_out_334( ArrayRowModule_2_io_V_wire_out_334 ),
       .io_V_wire_out_333( ArrayRowModule_2_io_V_wire_out_333 ),
       .io_V_wire_out_332( ArrayRowModule_2_io_V_wire_out_332 ),
       .io_V_wire_out_331( ArrayRowModule_2_io_V_wire_out_331 ),
       .io_V_wire_out_330( ArrayRowModule_2_io_V_wire_out_330 ),
       .io_V_wire_out_329( ArrayRowModule_2_io_V_wire_out_329 ),
       .io_V_wire_out_328( ArrayRowModule_2_io_V_wire_out_328 ),
       .io_V_wire_out_327( ArrayRowModule_2_io_V_wire_out_327 ),
       .io_V_wire_out_326( ArrayRowModule_2_io_V_wire_out_326 ),
       .io_V_wire_out_325( ArrayRowModule_2_io_V_wire_out_325 ),
       .io_V_wire_out_324( ArrayRowModule_2_io_V_wire_out_324 ),
       .io_V_wire_out_323( ArrayRowModule_2_io_V_wire_out_323 ),
       .io_V_wire_out_322( ArrayRowModule_2_io_V_wire_out_322 ),
       .io_V_wire_out_321( ArrayRowModule_2_io_V_wire_out_321 ),
       .io_V_wire_out_320( ArrayRowModule_2_io_V_wire_out_320 ),
       .io_V_wire_out_319( ArrayRowModule_2_io_V_wire_out_319 ),
       .io_V_wire_out_318( ArrayRowModule_2_io_V_wire_out_318 ),
       .io_V_wire_out_317( ArrayRowModule_2_io_V_wire_out_317 ),
       .io_V_wire_out_316( ArrayRowModule_2_io_V_wire_out_316 ),
       .io_V_wire_out_315( ArrayRowModule_2_io_V_wire_out_315 ),
       .io_V_wire_out_314( ArrayRowModule_2_io_V_wire_out_314 ),
       .io_V_wire_out_313( ArrayRowModule_2_io_V_wire_out_313 ),
       .io_V_wire_out_312( ArrayRowModule_2_io_V_wire_out_312 ),
       .io_V_wire_out_311( ArrayRowModule_2_io_V_wire_out_311 ),
       .io_V_wire_out_310( ArrayRowModule_2_io_V_wire_out_310 ),
       .io_V_wire_out_309( ArrayRowModule_2_io_V_wire_out_309 ),
       .io_V_wire_out_308( ArrayRowModule_2_io_V_wire_out_308 ),
       .io_V_wire_out_307( ArrayRowModule_2_io_V_wire_out_307 ),
       .io_V_wire_out_306( ArrayRowModule_2_io_V_wire_out_306 ),
       .io_V_wire_out_305( ArrayRowModule_2_io_V_wire_out_305 ),
       .io_V_wire_out_304( ArrayRowModule_2_io_V_wire_out_304 ),
       .io_V_wire_out_303( ArrayRowModule_2_io_V_wire_out_303 ),
       .io_V_wire_out_302( ArrayRowModule_2_io_V_wire_out_302 ),
       .io_V_wire_out_301( ArrayRowModule_2_io_V_wire_out_301 ),
       .io_V_wire_out_300( ArrayRowModule_2_io_V_wire_out_300 ),
       .io_V_wire_out_299( ArrayRowModule_2_io_V_wire_out_299 ),
       .io_V_wire_out_298( ArrayRowModule_2_io_V_wire_out_298 ),
       .io_V_wire_out_297( ArrayRowModule_2_io_V_wire_out_297 ),
       .io_V_wire_out_296( ArrayRowModule_2_io_V_wire_out_296 ),
       .io_V_wire_out_295( ArrayRowModule_2_io_V_wire_out_295 ),
       .io_V_wire_out_294( ArrayRowModule_2_io_V_wire_out_294 ),
       .io_V_wire_out_293( ArrayRowModule_2_io_V_wire_out_293 ),
       .io_V_wire_out_292( ArrayRowModule_2_io_V_wire_out_292 ),
       .io_V_wire_out_291( ArrayRowModule_2_io_V_wire_out_291 ),
       .io_V_wire_out_290( ArrayRowModule_2_io_V_wire_out_290 ),
       .io_V_wire_out_289( ArrayRowModule_2_io_V_wire_out_289 ),
       .io_V_wire_out_288( ArrayRowModule_2_io_V_wire_out_288 ),
       .io_V_wire_out_287( ArrayRowModule_2_io_V_wire_out_287 ),
       .io_V_wire_out_286( ArrayRowModule_2_io_V_wire_out_286 ),
       .io_V_wire_out_285( ArrayRowModule_2_io_V_wire_out_285 ),
       .io_V_wire_out_284( ArrayRowModule_2_io_V_wire_out_284 ),
       .io_V_wire_out_283( ArrayRowModule_2_io_V_wire_out_283 ),
       .io_V_wire_out_282( ArrayRowModule_2_io_V_wire_out_282 ),
       .io_V_wire_out_281( ArrayRowModule_2_io_V_wire_out_281 ),
       .io_V_wire_out_280( ArrayRowModule_2_io_V_wire_out_280 ),
       .io_V_wire_out_279( ArrayRowModule_2_io_V_wire_out_279 ),
       .io_V_wire_out_278( ArrayRowModule_2_io_V_wire_out_278 ),
       .io_V_wire_out_277( ArrayRowModule_2_io_V_wire_out_277 ),
       .io_V_wire_out_276( ArrayRowModule_2_io_V_wire_out_276 ),
       .io_V_wire_out_275( ArrayRowModule_2_io_V_wire_out_275 ),
       .io_V_wire_out_274( ArrayRowModule_2_io_V_wire_out_274 ),
       .io_V_wire_out_273( ArrayRowModule_2_io_V_wire_out_273 ),
       .io_V_wire_out_272( ArrayRowModule_2_io_V_wire_out_272 ),
       .io_V_wire_out_271( ArrayRowModule_2_io_V_wire_out_271 ),
       .io_V_wire_out_270( ArrayRowModule_2_io_V_wire_out_270 ),
       .io_V_wire_out_269( ArrayRowModule_2_io_V_wire_out_269 ),
       .io_V_wire_out_268( ArrayRowModule_2_io_V_wire_out_268 ),
       .io_V_wire_out_267( ArrayRowModule_2_io_V_wire_out_267 ),
       .io_V_wire_out_266( ArrayRowModule_2_io_V_wire_out_266 ),
       .io_V_wire_out_265( ArrayRowModule_2_io_V_wire_out_265 ),
       .io_V_wire_out_264( ArrayRowModule_2_io_V_wire_out_264 ),
       .io_V_wire_out_263( ArrayRowModule_2_io_V_wire_out_263 ),
       .io_V_wire_out_262( ArrayRowModule_2_io_V_wire_out_262 ),
       .io_V_wire_out_261( ArrayRowModule_2_io_V_wire_out_261 ),
       .io_V_wire_out_260( ArrayRowModule_2_io_V_wire_out_260 ),
       .io_V_wire_out_259( ArrayRowModule_2_io_V_wire_out_259 ),
       .io_V_wire_out_258( ArrayRowModule_2_io_V_wire_out_258 ),
       .io_V_wire_out_257( ArrayRowModule_2_io_V_wire_out_257 ),
       .io_V_wire_out_256( ArrayRowModule_2_io_V_wire_out_256 ),
       .io_V_wire_out_255( ArrayRowModule_2_io_V_wire_out_255 ),
       .io_V_wire_out_254( ArrayRowModule_2_io_V_wire_out_254 ),
       .io_V_wire_out_253( ArrayRowModule_2_io_V_wire_out_253 ),
       .io_V_wire_out_252( ArrayRowModule_2_io_V_wire_out_252 ),
       .io_V_wire_out_251( ArrayRowModule_2_io_V_wire_out_251 ),
       .io_V_wire_out_250( ArrayRowModule_2_io_V_wire_out_250 ),
       .io_V_wire_out_249( ArrayRowModule_2_io_V_wire_out_249 ),
       .io_V_wire_out_248( ArrayRowModule_2_io_V_wire_out_248 ),
       .io_V_wire_out_247( ArrayRowModule_2_io_V_wire_out_247 ),
       .io_V_wire_out_246( ArrayRowModule_2_io_V_wire_out_246 ),
       .io_V_wire_out_245( ArrayRowModule_2_io_V_wire_out_245 ),
       .io_V_wire_out_244( ArrayRowModule_2_io_V_wire_out_244 ),
       .io_V_wire_out_243( ArrayRowModule_2_io_V_wire_out_243 ),
       .io_V_wire_out_242( ArrayRowModule_2_io_V_wire_out_242 ),
       .io_V_wire_out_241( ArrayRowModule_2_io_V_wire_out_241 ),
       .io_V_wire_out_240( ArrayRowModule_2_io_V_wire_out_240 ),
       .io_V_wire_out_239( ArrayRowModule_2_io_V_wire_out_239 ),
       .io_V_wire_out_238( ArrayRowModule_2_io_V_wire_out_238 ),
       .io_V_wire_out_237( ArrayRowModule_2_io_V_wire_out_237 ),
       .io_V_wire_out_236( ArrayRowModule_2_io_V_wire_out_236 ),
       .io_V_wire_out_235( ArrayRowModule_2_io_V_wire_out_235 ),
       .io_V_wire_out_234( ArrayRowModule_2_io_V_wire_out_234 ),
       .io_V_wire_out_233( ArrayRowModule_2_io_V_wire_out_233 ),
       .io_V_wire_out_232( ArrayRowModule_2_io_V_wire_out_232 ),
       .io_V_wire_out_231( ArrayRowModule_2_io_V_wire_out_231 ),
       .io_V_wire_out_230( ArrayRowModule_2_io_V_wire_out_230 ),
       .io_V_wire_out_229( ArrayRowModule_2_io_V_wire_out_229 ),
       .io_V_wire_out_228( ArrayRowModule_2_io_V_wire_out_228 ),
       .io_V_wire_out_227( ArrayRowModule_2_io_V_wire_out_227 ),
       .io_V_wire_out_226( ArrayRowModule_2_io_V_wire_out_226 ),
       .io_V_wire_out_225( ArrayRowModule_2_io_V_wire_out_225 ),
       .io_V_wire_out_224( ArrayRowModule_2_io_V_wire_out_224 ),
       .io_V_wire_out_223( ArrayRowModule_2_io_V_wire_out_223 ),
       .io_V_wire_out_222( ArrayRowModule_2_io_V_wire_out_222 ),
       .io_V_wire_out_221( ArrayRowModule_2_io_V_wire_out_221 ),
       .io_V_wire_out_220( ArrayRowModule_2_io_V_wire_out_220 ),
       .io_V_wire_out_219( ArrayRowModule_2_io_V_wire_out_219 ),
       .io_V_wire_out_218( ArrayRowModule_2_io_V_wire_out_218 ),
       .io_V_wire_out_217( ArrayRowModule_2_io_V_wire_out_217 ),
       .io_V_wire_out_216( ArrayRowModule_2_io_V_wire_out_216 ),
       .io_V_wire_out_215( ArrayRowModule_2_io_V_wire_out_215 ),
       .io_V_wire_out_214( ArrayRowModule_2_io_V_wire_out_214 ),
       .io_V_wire_out_213( ArrayRowModule_2_io_V_wire_out_213 ),
       .io_V_wire_out_212( ArrayRowModule_2_io_V_wire_out_212 ),
       .io_V_wire_out_211( ArrayRowModule_2_io_V_wire_out_211 ),
       .io_V_wire_out_210( ArrayRowModule_2_io_V_wire_out_210 ),
       .io_V_wire_out_209( ArrayRowModule_2_io_V_wire_out_209 ),
       .io_V_wire_out_208( ArrayRowModule_2_io_V_wire_out_208 ),
       .io_V_wire_out_207( ArrayRowModule_2_io_V_wire_out_207 ),
       .io_V_wire_out_206( ArrayRowModule_2_io_V_wire_out_206 ),
       .io_V_wire_out_205( ArrayRowModule_2_io_V_wire_out_205 ),
       .io_V_wire_out_204( ArrayRowModule_2_io_V_wire_out_204 ),
       .io_V_wire_out_203( ArrayRowModule_2_io_V_wire_out_203 ),
       .io_V_wire_out_202( ArrayRowModule_2_io_V_wire_out_202 ),
       .io_V_wire_out_201( ArrayRowModule_2_io_V_wire_out_201 ),
       .io_V_wire_out_200( ArrayRowModule_2_io_V_wire_out_200 ),
       .io_V_wire_out_199( ArrayRowModule_2_io_V_wire_out_199 ),
       .io_V_wire_out_198( ArrayRowModule_2_io_V_wire_out_198 ),
       .io_V_wire_out_197( ArrayRowModule_2_io_V_wire_out_197 ),
       .io_V_wire_out_196( ArrayRowModule_2_io_V_wire_out_196 ),
       .io_V_wire_out_195( ArrayRowModule_2_io_V_wire_out_195 ),
       .io_V_wire_out_194( ArrayRowModule_2_io_V_wire_out_194 ),
       .io_V_wire_out_193( ArrayRowModule_2_io_V_wire_out_193 ),
       .io_V_wire_out_192( ArrayRowModule_2_io_V_wire_out_192 ),
       .io_V_wire_out_191( ArrayRowModule_2_io_V_wire_out_191 ),
       .io_V_wire_out_190( ArrayRowModule_2_io_V_wire_out_190 ),
       .io_V_wire_out_189( ArrayRowModule_2_io_V_wire_out_189 ),
       .io_V_wire_out_188( ArrayRowModule_2_io_V_wire_out_188 ),
       .io_V_wire_out_187( ArrayRowModule_2_io_V_wire_out_187 ),
       .io_V_wire_out_186( ArrayRowModule_2_io_V_wire_out_186 ),
       .io_V_wire_out_185( ArrayRowModule_2_io_V_wire_out_185 ),
       .io_V_wire_out_184( ArrayRowModule_2_io_V_wire_out_184 ),
       .io_V_wire_out_183( ArrayRowModule_2_io_V_wire_out_183 ),
       .io_V_wire_out_182( ArrayRowModule_2_io_V_wire_out_182 ),
       .io_V_wire_out_181( ArrayRowModule_2_io_V_wire_out_181 ),
       .io_V_wire_out_180( ArrayRowModule_2_io_V_wire_out_180 ),
       .io_V_wire_out_179( ArrayRowModule_2_io_V_wire_out_179 ),
       .io_V_wire_out_178( ArrayRowModule_2_io_V_wire_out_178 ),
       .io_V_wire_out_177( ArrayRowModule_2_io_V_wire_out_177 ),
       .io_V_wire_out_176( ArrayRowModule_2_io_V_wire_out_176 ),
       .io_V_wire_out_175( ArrayRowModule_2_io_V_wire_out_175 ),
       .io_V_wire_out_174( ArrayRowModule_2_io_V_wire_out_174 ),
       .io_V_wire_out_173( ArrayRowModule_2_io_V_wire_out_173 ),
       .io_V_wire_out_172( ArrayRowModule_2_io_V_wire_out_172 ),
       .io_V_wire_out_171( ArrayRowModule_2_io_V_wire_out_171 ),
       .io_V_wire_out_170( ArrayRowModule_2_io_V_wire_out_170 ),
       .io_V_wire_out_169( ArrayRowModule_2_io_V_wire_out_169 ),
       .io_V_wire_out_168( ArrayRowModule_2_io_V_wire_out_168 ),
       .io_V_wire_out_167( ArrayRowModule_2_io_V_wire_out_167 ),
       .io_V_wire_out_166( ArrayRowModule_2_io_V_wire_out_166 ),
       .io_V_wire_out_165( ArrayRowModule_2_io_V_wire_out_165 ),
       .io_V_wire_out_164( ArrayRowModule_2_io_V_wire_out_164 ),
       .io_V_wire_out_163( ArrayRowModule_2_io_V_wire_out_163 ),
       .io_V_wire_out_162( ArrayRowModule_2_io_V_wire_out_162 ),
       .io_V_wire_out_161( ArrayRowModule_2_io_V_wire_out_161 ),
       .io_V_wire_out_160( ArrayRowModule_2_io_V_wire_out_160 ),
       .io_V_wire_out_159( ArrayRowModule_2_io_V_wire_out_159 ),
       .io_V_wire_out_158( ArrayRowModule_2_io_V_wire_out_158 ),
       .io_V_wire_out_157( ArrayRowModule_2_io_V_wire_out_157 ),
       .io_V_wire_out_156( ArrayRowModule_2_io_V_wire_out_156 ),
       .io_V_wire_out_155( ArrayRowModule_2_io_V_wire_out_155 ),
       .io_V_wire_out_154( ArrayRowModule_2_io_V_wire_out_154 ),
       .io_V_wire_out_153( ArrayRowModule_2_io_V_wire_out_153 ),
       .io_V_wire_out_152( ArrayRowModule_2_io_V_wire_out_152 ),
       .io_V_wire_out_151( ArrayRowModule_2_io_V_wire_out_151 ),
       .io_V_wire_out_150( ArrayRowModule_2_io_V_wire_out_150 ),
       .io_V_wire_out_149( ArrayRowModule_2_io_V_wire_out_149 ),
       .io_V_wire_out_148( ArrayRowModule_2_io_V_wire_out_148 ),
       .io_V_wire_out_147( ArrayRowModule_2_io_V_wire_out_147 ),
       .io_V_wire_out_146( ArrayRowModule_2_io_V_wire_out_146 ),
       .io_V_wire_out_145( ArrayRowModule_2_io_V_wire_out_145 ),
       .io_V_wire_out_144( ArrayRowModule_2_io_V_wire_out_144 ),
       .io_V_wire_out_143( ArrayRowModule_2_io_V_wire_out_143 ),
       .io_V_wire_out_142( ArrayRowModule_2_io_V_wire_out_142 ),
       .io_V_wire_out_141( ArrayRowModule_2_io_V_wire_out_141 ),
       .io_V_wire_out_140( ArrayRowModule_2_io_V_wire_out_140 ),
       .io_V_wire_out_139( ArrayRowModule_2_io_V_wire_out_139 ),
       .io_V_wire_out_138( ArrayRowModule_2_io_V_wire_out_138 ),
       .io_V_wire_out_137( ArrayRowModule_2_io_V_wire_out_137 ),
       .io_V_wire_out_136( ArrayRowModule_2_io_V_wire_out_136 ),
       .io_V_wire_out_135( ArrayRowModule_2_io_V_wire_out_135 ),
       .io_V_wire_out_134( ArrayRowModule_2_io_V_wire_out_134 ),
       .io_V_wire_out_133( ArrayRowModule_2_io_V_wire_out_133 ),
       .io_V_wire_out_132( ArrayRowModule_2_io_V_wire_out_132 ),
       .io_V_wire_out_131( ArrayRowModule_2_io_V_wire_out_131 ),
       .io_V_wire_out_130( ArrayRowModule_2_io_V_wire_out_130 ),
       .io_V_wire_out_129( ArrayRowModule_2_io_V_wire_out_129 ),
       .io_V_wire_out_128( ArrayRowModule_2_io_V_wire_out_128 ),
       .io_V_wire_out_127( ArrayRowModule_2_io_V_wire_out_127 ),
       .io_V_wire_out_126( ArrayRowModule_2_io_V_wire_out_126 ),
       .io_V_wire_out_125( ArrayRowModule_2_io_V_wire_out_125 ),
       .io_V_wire_out_124( ArrayRowModule_2_io_V_wire_out_124 ),
       .io_V_wire_out_123( ArrayRowModule_2_io_V_wire_out_123 ),
       .io_V_wire_out_122( ArrayRowModule_2_io_V_wire_out_122 ),
       .io_V_wire_out_121( ArrayRowModule_2_io_V_wire_out_121 ),
       .io_V_wire_out_120( ArrayRowModule_2_io_V_wire_out_120 ),
       .io_V_wire_out_119( ArrayRowModule_2_io_V_wire_out_119 ),
       .io_V_wire_out_118( ArrayRowModule_2_io_V_wire_out_118 ),
       .io_V_wire_out_117( ArrayRowModule_2_io_V_wire_out_117 ),
       .io_V_wire_out_116( ArrayRowModule_2_io_V_wire_out_116 ),
       .io_V_wire_out_115( ArrayRowModule_2_io_V_wire_out_115 ),
       .io_V_wire_out_114( ArrayRowModule_2_io_V_wire_out_114 ),
       .io_V_wire_out_113( ArrayRowModule_2_io_V_wire_out_113 ),
       .io_V_wire_out_112( ArrayRowModule_2_io_V_wire_out_112 ),
       .io_V_wire_out_111( ArrayRowModule_2_io_V_wire_out_111 ),
       .io_V_wire_out_110( ArrayRowModule_2_io_V_wire_out_110 ),
       .io_V_wire_out_109( ArrayRowModule_2_io_V_wire_out_109 ),
       .io_V_wire_out_108( ArrayRowModule_2_io_V_wire_out_108 ),
       .io_V_wire_out_107( ArrayRowModule_2_io_V_wire_out_107 ),
       .io_V_wire_out_106( ArrayRowModule_2_io_V_wire_out_106 ),
       .io_V_wire_out_105( ArrayRowModule_2_io_V_wire_out_105 ),
       .io_V_wire_out_104( ArrayRowModule_2_io_V_wire_out_104 ),
       .io_V_wire_out_103( ArrayRowModule_2_io_V_wire_out_103 ),
       .io_V_wire_out_102( ArrayRowModule_2_io_V_wire_out_102 ),
       .io_V_wire_out_101( ArrayRowModule_2_io_V_wire_out_101 ),
       .io_V_wire_out_100( ArrayRowModule_2_io_V_wire_out_100 ),
       .io_V_wire_out_99( ArrayRowModule_2_io_V_wire_out_99 ),
       .io_V_wire_out_98( ArrayRowModule_2_io_V_wire_out_98 ),
       .io_V_wire_out_97( ArrayRowModule_2_io_V_wire_out_97 ),
       .io_V_wire_out_96( ArrayRowModule_2_io_V_wire_out_96 ),
       .io_V_wire_out_95( ArrayRowModule_2_io_V_wire_out_95 ),
       .io_V_wire_out_94( ArrayRowModule_2_io_V_wire_out_94 ),
       .io_V_wire_out_93( ArrayRowModule_2_io_V_wire_out_93 ),
       .io_V_wire_out_92( ArrayRowModule_2_io_V_wire_out_92 ),
       .io_V_wire_out_91( ArrayRowModule_2_io_V_wire_out_91 ),
       .io_V_wire_out_90( ArrayRowModule_2_io_V_wire_out_90 ),
       .io_V_wire_out_89( ArrayRowModule_2_io_V_wire_out_89 ),
       .io_V_wire_out_88( ArrayRowModule_2_io_V_wire_out_88 ),
       .io_V_wire_out_87( ArrayRowModule_2_io_V_wire_out_87 ),
       .io_V_wire_out_86( ArrayRowModule_2_io_V_wire_out_86 ),
       .io_V_wire_out_85( ArrayRowModule_2_io_V_wire_out_85 ),
       .io_V_wire_out_84( ArrayRowModule_2_io_V_wire_out_84 ),
       .io_V_wire_out_83( ArrayRowModule_2_io_V_wire_out_83 ),
       .io_V_wire_out_82( ArrayRowModule_2_io_V_wire_out_82 ),
       .io_V_wire_out_81( ArrayRowModule_2_io_V_wire_out_81 ),
       .io_V_wire_out_80( ArrayRowModule_2_io_V_wire_out_80 ),
       .io_V_wire_out_79( ArrayRowModule_2_io_V_wire_out_79 ),
       .io_V_wire_out_78( ArrayRowModule_2_io_V_wire_out_78 ),
       .io_V_wire_out_77( ArrayRowModule_2_io_V_wire_out_77 ),
       .io_V_wire_out_76( ArrayRowModule_2_io_V_wire_out_76 ),
       .io_V_wire_out_75( ArrayRowModule_2_io_V_wire_out_75 ),
       .io_V_wire_out_74( ArrayRowModule_2_io_V_wire_out_74 ),
       .io_V_wire_out_73( ArrayRowModule_2_io_V_wire_out_73 ),
       .io_V_wire_out_72( ArrayRowModule_2_io_V_wire_out_72 ),
       .io_V_wire_out_71( ArrayRowModule_2_io_V_wire_out_71 ),
       .io_V_wire_out_70( ArrayRowModule_2_io_V_wire_out_70 ),
       .io_V_wire_out_69( ArrayRowModule_2_io_V_wire_out_69 ),
       .io_V_wire_out_68( ArrayRowModule_2_io_V_wire_out_68 ),
       .io_V_wire_out_67( ArrayRowModule_2_io_V_wire_out_67 ),
       .io_V_wire_out_66( ArrayRowModule_2_io_V_wire_out_66 ),
       .io_V_wire_out_65( ArrayRowModule_2_io_V_wire_out_65 ),
       .io_V_wire_out_64( ArrayRowModule_2_io_V_wire_out_64 ),
       .io_V_wire_out_63( ArrayRowModule_2_io_V_wire_out_63 ),
       .io_V_wire_out_62( ArrayRowModule_2_io_V_wire_out_62 ),
       .io_V_wire_out_61( ArrayRowModule_2_io_V_wire_out_61 ),
       .io_V_wire_out_60( ArrayRowModule_2_io_V_wire_out_60 ),
       .io_V_wire_out_59( ArrayRowModule_2_io_V_wire_out_59 ),
       .io_V_wire_out_58( ArrayRowModule_2_io_V_wire_out_58 ),
       .io_V_wire_out_57( ArrayRowModule_2_io_V_wire_out_57 ),
       .io_V_wire_out_56( ArrayRowModule_2_io_V_wire_out_56 ),
       .io_V_wire_out_55( ArrayRowModule_2_io_V_wire_out_55 ),
       .io_V_wire_out_54( ArrayRowModule_2_io_V_wire_out_54 ),
       .io_V_wire_out_53( ArrayRowModule_2_io_V_wire_out_53 ),
       .io_V_wire_out_52( ArrayRowModule_2_io_V_wire_out_52 ),
       .io_V_wire_out_51( ArrayRowModule_2_io_V_wire_out_51 ),
       .io_V_wire_out_50( ArrayRowModule_2_io_V_wire_out_50 ),
       .io_V_wire_out_49( ArrayRowModule_2_io_V_wire_out_49 ),
       .io_V_wire_out_48( ArrayRowModule_2_io_V_wire_out_48 ),
       .io_V_wire_out_47( ArrayRowModule_2_io_V_wire_out_47 ),
       .io_V_wire_out_46( ArrayRowModule_2_io_V_wire_out_46 ),
       .io_V_wire_out_45( ArrayRowModule_2_io_V_wire_out_45 ),
       .io_V_wire_out_44( ArrayRowModule_2_io_V_wire_out_44 ),
       .io_V_wire_out_43( ArrayRowModule_2_io_V_wire_out_43 ),
       .io_V_wire_out_42( ArrayRowModule_2_io_V_wire_out_42 ),
       .io_V_wire_out_41( ArrayRowModule_2_io_V_wire_out_41 ),
       .io_V_wire_out_40( ArrayRowModule_2_io_V_wire_out_40 ),
       .io_V_wire_out_39( ArrayRowModule_2_io_V_wire_out_39 ),
       .io_V_wire_out_38( ArrayRowModule_2_io_V_wire_out_38 ),
       .io_V_wire_out_37( ArrayRowModule_2_io_V_wire_out_37 ),
       .io_V_wire_out_36( ArrayRowModule_2_io_V_wire_out_36 ),
       .io_V_wire_out_35( ArrayRowModule_2_io_V_wire_out_35 ),
       .io_V_wire_out_34( ArrayRowModule_2_io_V_wire_out_34 ),
       .io_V_wire_out_33( ArrayRowModule_2_io_V_wire_out_33 ),
       .io_V_wire_out_32( ArrayRowModule_2_io_V_wire_out_32 ),
       .io_V_wire_out_31( ArrayRowModule_2_io_V_wire_out_31 ),
       .io_V_wire_out_30( ArrayRowModule_2_io_V_wire_out_30 ),
       .io_V_wire_out_29( ArrayRowModule_2_io_V_wire_out_29 ),
       .io_V_wire_out_28( ArrayRowModule_2_io_V_wire_out_28 ),
       .io_V_wire_out_27( ArrayRowModule_2_io_V_wire_out_27 ),
       .io_V_wire_out_26( ArrayRowModule_2_io_V_wire_out_26 ),
       .io_V_wire_out_25( ArrayRowModule_2_io_V_wire_out_25 ),
       .io_V_wire_out_24( ArrayRowModule_2_io_V_wire_out_24 ),
       .io_V_wire_out_23( ArrayRowModule_2_io_V_wire_out_23 ),
       .io_V_wire_out_22( ArrayRowModule_2_io_V_wire_out_22 ),
       .io_V_wire_out_21( ArrayRowModule_2_io_V_wire_out_21 ),
       .io_V_wire_out_20( ArrayRowModule_2_io_V_wire_out_20 ),
       .io_V_wire_out_19( ArrayRowModule_2_io_V_wire_out_19 ),
       .io_V_wire_out_18( ArrayRowModule_2_io_V_wire_out_18 ),
       .io_V_wire_out_17( ArrayRowModule_2_io_V_wire_out_17 ),
       .io_V_wire_out_16( ArrayRowModule_2_io_V_wire_out_16 ),
       .io_V_wire_out_15( ArrayRowModule_2_io_V_wire_out_15 ),
       .io_V_wire_out_14( ArrayRowModule_2_io_V_wire_out_14 ),
       .io_V_wire_out_13( ArrayRowModule_2_io_V_wire_out_13 ),
       .io_V_wire_out_12( ArrayRowModule_2_io_V_wire_out_12 ),
       .io_V_wire_out_11( ArrayRowModule_2_io_V_wire_out_11 ),
       .io_V_wire_out_10( ArrayRowModule_2_io_V_wire_out_10 ),
       .io_V_wire_out_9( ArrayRowModule_2_io_V_wire_out_9 ),
       .io_V_wire_out_8( ArrayRowModule_2_io_V_wire_out_8 ),
       .io_V_wire_out_7( ArrayRowModule_2_io_V_wire_out_7 ),
       .io_V_wire_out_6( ArrayRowModule_2_io_V_wire_out_6 ),
       .io_V_wire_out_5( ArrayRowModule_2_io_V_wire_out_5 ),
       .io_V_wire_out_4( ArrayRowModule_2_io_V_wire_out_4 ),
       .io_V_wire_out_3( ArrayRowModule_2_io_V_wire_out_3 ),
       .io_V_wire_out_2( ArrayRowModule_2_io_V_wire_out_2 ),
       .io_V_wire_out_1( ArrayRowModule_2_io_V_wire_out_1 ),
       .io_V_wire_out_0( ArrayRowModule_2_io_V_wire_out_0 ),
       .io_V_wire_en_22( ArrayRowModule_2_io_V_wire_en_22 ),
       .io_V_wire_en_21( ArrayRowModule_2_io_V_wire_en_21 ),
       .io_V_wire_en_20( ArrayRowModule_2_io_V_wire_en_20 ),
       .io_V_wire_en_19( ArrayRowModule_2_io_V_wire_en_19 ),
       .io_V_wire_en_18( ArrayRowModule_2_io_V_wire_en_18 ),
       .io_V_wire_en_17( ArrayRowModule_2_io_V_wire_en_17 ),
       .io_V_wire_en_16( ArrayRowModule_2_io_V_wire_en_16 ),
       .io_V_wire_en_15( ArrayRowModule_2_io_V_wire_en_15 ),
       .io_V_wire_en_14( ArrayRowModule_2_io_V_wire_en_14 ),
       .io_V_wire_en_13( ArrayRowModule_2_io_V_wire_en_13 ),
       .io_V_wire_en_12( ArrayRowModule_2_io_V_wire_en_12 ),
       .io_V_wire_en_11( ArrayRowModule_2_io_V_wire_en_11 ),
       .io_V_wire_en_10( ArrayRowModule_2_io_V_wire_en_10 ),
       .io_V_wire_en_9( ArrayRowModule_2_io_V_wire_en_9 ),
       .io_V_wire_en_8( ArrayRowModule_2_io_V_wire_en_8 ),
       .io_V_wire_en_7( ArrayRowModule_2_io_V_wire_en_7 ),
       .io_V_wire_en_6( ArrayRowModule_2_io_V_wire_en_6 ),
       .io_V_wire_en_5( ArrayRowModule_2_io_V_wire_en_5 ),
       .io_V_wire_en_4( ArrayRowModule_2_io_V_wire_en_4 ),
       .io_V_wire_en_3( ArrayRowModule_2_io_V_wire_en_3 ),
       .io_V_wire_en_2( ArrayRowModule_2_io_V_wire_en_2 ),
       .io_V_wire_en_1( ArrayRowModule_2_io_V_wire_en_1 ),
       .io_V_wire_en_0( ArrayRowModule_2_io_V_wire_en_0 ),
       .io_G_wire_above_3( ArrayRowModule_1_io_G_wire_below_3 ),
       .io_G_wire_above_2( ArrayRowModule_1_io_G_wire_below_2 ),
       .io_G_wire_above_1( ArrayRowModule_1_io_G_wire_below_1 ),
       .io_G_wire_above_0( ArrayRowModule_1_io_G_wire_below_0 ),
       .io_H_wire_above_32( ArrayRowModule_1_io_H_wire_below_32 ),
       .io_H_wire_above_31( ArrayRowModule_1_io_H_wire_below_31 ),
       .io_H_wire_above_30( ArrayRowModule_1_io_H_wire_below_30 ),
       .io_H_wire_above_29( ArrayRowModule_1_io_H_wire_below_29 ),
       .io_H_wire_above_28( ArrayRowModule_1_io_H_wire_below_28 ),
       .io_H_wire_above_27( ArrayRowModule_1_io_H_wire_below_27 ),
       .io_H_wire_above_26( ArrayRowModule_1_io_H_wire_below_26 ),
       .io_H_wire_above_25( ArrayRowModule_1_io_H_wire_below_25 ),
       .io_H_wire_above_24( ArrayRowModule_1_io_H_wire_below_24 ),
       .io_H_wire_above_23( ArrayRowModule_1_io_H_wire_below_23 ),
       .io_H_wire_above_22( ArrayRowModule_1_io_H_wire_below_22 ),
       .io_H_wire_above_21( ArrayRowModule_1_io_H_wire_below_21 ),
       .io_H_wire_above_20( ArrayRowModule_1_io_H_wire_below_20 ),
       .io_H_wire_above_19( ArrayRowModule_1_io_H_wire_below_19 ),
       .io_H_wire_above_18( ArrayRowModule_1_io_H_wire_below_18 ),
       .io_H_wire_above_17( ArrayRowModule_1_io_H_wire_below_17 ),
       .io_H_wire_above_16( ArrayRowModule_1_io_H_wire_below_16 ),
       .io_H_wire_above_15( ArrayRowModule_1_io_H_wire_below_15 ),
       .io_H_wire_above_14( ArrayRowModule_1_io_H_wire_below_14 ),
       .io_H_wire_above_13( ArrayRowModule_1_io_H_wire_below_13 ),
       .io_H_wire_above_12( ArrayRowModule_1_io_H_wire_below_12 ),
       .io_H_wire_above_11( ArrayRowModule_1_io_H_wire_below_11 ),
       .io_H_wire_above_10( ArrayRowModule_1_io_H_wire_below_10 ),
       .io_H_wire_above_9( ArrayRowModule_1_io_H_wire_below_9 ),
       .io_H_wire_above_8( ArrayRowModule_1_io_H_wire_below_8 ),
       .io_H_wire_above_7( ArrayRowModule_1_io_H_wire_below_7 ),
       .io_H_wire_above_6( ArrayRowModule_1_io_H_wire_below_6 ),
       .io_H_wire_above_5( ArrayRowModule_1_io_H_wire_below_5 ),
       .io_H_wire_above_4( ArrayRowModule_1_io_H_wire_below_4 ),
       .io_H_wire_above_3( ArrayRowModule_1_io_H_wire_below_3 ),
       .io_H_wire_above_2( ArrayRowModule_1_io_H_wire_below_2 ),
       .io_H_wire_above_1( ArrayRowModule_1_io_H_wire_below_1 ),
       .io_H_wire_above_0( ArrayRowModule_1_io_H_wire_below_0 ),
       .io_mem_bus_in_23( ArrayRowModule_1_io_mem_bus_out_23 ),
       .io_mem_bus_in_22( ArrayRowModule_1_io_mem_bus_out_22 ),
       .io_mem_bus_in_21( ArrayRowModule_1_io_mem_bus_out_21 ),
       .io_mem_bus_in_20( ArrayRowModule_1_io_mem_bus_out_20 ),
       .io_mem_bus_in_19( ArrayRowModule_1_io_mem_bus_out_19 ),
       .io_mem_bus_in_18( ArrayRowModule_1_io_mem_bus_out_18 ),
       .io_mem_bus_in_17( ArrayRowModule_1_io_mem_bus_out_17 ),
       .io_mem_bus_in_16( ArrayRowModule_1_io_mem_bus_out_16 ),
       .io_mem_bus_in_15( ArrayRowModule_1_io_mem_bus_out_15 ),
       .io_mem_bus_in_14( ArrayRowModule_1_io_mem_bus_out_14 ),
       .io_mem_bus_in_13( ArrayRowModule_1_io_mem_bus_out_13 ),
       .io_mem_bus_in_12( ArrayRowModule_1_io_mem_bus_out_12 ),
       .io_mem_bus_in_11( ArrayRowModule_1_io_mem_bus_out_11 ),
       .io_mem_bus_in_10( ArrayRowModule_1_io_mem_bus_out_10 ),
       .io_mem_bus_in_9( ArrayRowModule_1_io_mem_bus_out_9 ),
       .io_mem_bus_in_8( ArrayRowModule_1_io_mem_bus_out_8 ),
       .io_mem_bus_in_7( ArrayRowModule_1_io_mem_bus_out_7 ),
       .io_mem_bus_in_6( ArrayRowModule_1_io_mem_bus_out_6 ),
       .io_mem_bus_in_5( ArrayRowModule_1_io_mem_bus_out_5 ),
       .io_mem_bus_in_4( ArrayRowModule_1_io_mem_bus_out_4 ),
       .io_mem_bus_in_3( ArrayRowModule_1_io_mem_bus_out_3 ),
       .io_mem_bus_in_2( ArrayRowModule_1_io_mem_bus_out_2 ),
       .io_mem_bus_in_1( ArrayRowModule_1_io_mem_bus_out_1 ),
       .io_mem_bus_in_0( ArrayRowModule_1_io_mem_bus_out_0 ),
       .io_H_out_above_22( ArrayRowModule_1_io_H_out_22 ),
       .io_H_out_above_21( ArrayRowModule_1_io_H_out_21 ),
       .io_H_out_above_20( ArrayRowModule_1_io_H_out_20 ),
       .io_H_out_above_19( ArrayRowModule_1_io_H_out_19 ),
       .io_H_out_above_18( ArrayRowModule_1_io_H_out_18 ),
       .io_H_out_above_17( ArrayRowModule_1_io_H_out_17 ),
       .io_H_out_above_16( ArrayRowModule_1_io_H_out_16 ),
       .io_H_out_above_15( ArrayRowModule_1_io_H_out_15 ),
       .io_H_out_above_14( ArrayRowModule_1_io_H_out_14 ),
       .io_H_out_above_13( ArrayRowModule_1_io_H_out_13 ),
       .io_H_out_above_12( ArrayRowModule_1_io_H_out_12 ),
       .io_H_out_above_11( ArrayRowModule_1_io_H_out_11 ),
       .io_H_out_above_10( ArrayRowModule_1_io_H_out_10 ),
       .io_H_out_above_9( ArrayRowModule_1_io_H_out_9 ),
       .io_H_out_above_8( ArrayRowModule_1_io_H_out_8 ),
       .io_H_out_above_7( ArrayRowModule_1_io_H_out_7 ),
       .io_H_out_above_6( ArrayRowModule_1_io_H_out_6 ),
       .io_H_out_above_5( ArrayRowModule_1_io_H_out_5 ),
       .io_H_out_above_4( ArrayRowModule_1_io_H_out_4 ),
       .io_H_out_above_3( ArrayRowModule_1_io_H_out_3 ),
       .io_H_out_above_2( ArrayRowModule_1_io_H_out_2 ),
       .io_H_out_above_1( ArrayRowModule_1_io_H_out_1 ),
       .io_H_out_above_0( ArrayRowModule_1_io_H_out_0 ),
       .io_H_out_22( ArrayRowModule_2_io_H_out_22 ),
       .io_H_out_21( ArrayRowModule_2_io_H_out_21 ),
       .io_H_out_20( ArrayRowModule_2_io_H_out_20 ),
       .io_H_out_19( ArrayRowModule_2_io_H_out_19 ),
       .io_H_out_18( ArrayRowModule_2_io_H_out_18 ),
       .io_H_out_17( ArrayRowModule_2_io_H_out_17 ),
       .io_H_out_16( ArrayRowModule_2_io_H_out_16 ),
       .io_H_out_15( ArrayRowModule_2_io_H_out_15 ),
       .io_H_out_14( ArrayRowModule_2_io_H_out_14 ),
       .io_H_out_13( ArrayRowModule_2_io_H_out_13 ),
       .io_H_out_12( ArrayRowModule_2_io_H_out_12 ),
       .io_H_out_11( ArrayRowModule_2_io_H_out_11 ),
       .io_H_out_10( ArrayRowModule_2_io_H_out_10 ),
       .io_H_out_9( ArrayRowModule_2_io_H_out_9 ),
       .io_H_out_8( ArrayRowModule_2_io_H_out_8 ),
       .io_H_out_7( ArrayRowModule_2_io_H_out_7 ),
       .io_H_out_6( ArrayRowModule_2_io_H_out_6 ),
       .io_H_out_5( ArrayRowModule_2_io_H_out_5 ),
       .io_H_out_4( ArrayRowModule_2_io_H_out_4 ),
       .io_H_out_3( ArrayRowModule_2_io_H_out_3 ),
       .io_H_out_2( ArrayRowModule_2_io_H_out_2 ),
       .io_H_out_1( ArrayRowModule_2_io_H_out_1 ),
       .io_H_out_0( ArrayRowModule_2_io_H_out_0 ),
       .io_G_wire_below_3( ArrayRowModule_2_io_G_wire_below_3 ),
       .io_G_wire_below_2( ArrayRowModule_2_io_G_wire_below_2 ),
       .io_G_wire_below_1( ArrayRowModule_2_io_G_wire_below_1 ),
       .io_G_wire_below_0( ArrayRowModule_2_io_G_wire_below_0 ),
       .io_H_wire_below_32( ArrayRowModule_2_io_H_wire_below_32 ),
       .io_H_wire_below_31( ArrayRowModule_2_io_H_wire_below_31 ),
       .io_H_wire_below_30( ArrayRowModule_2_io_H_wire_below_30 ),
       .io_H_wire_below_29( ArrayRowModule_2_io_H_wire_below_29 ),
       .io_H_wire_below_28( ArrayRowModule_2_io_H_wire_below_28 ),
       .io_H_wire_below_27( ArrayRowModule_2_io_H_wire_below_27 ),
       .io_H_wire_below_26( ArrayRowModule_2_io_H_wire_below_26 ),
       .io_H_wire_below_25( ArrayRowModule_2_io_H_wire_below_25 ),
       .io_H_wire_below_24( ArrayRowModule_2_io_H_wire_below_24 ),
       .io_H_wire_below_23( ArrayRowModule_2_io_H_wire_below_23 ),
       .io_H_wire_below_22( ArrayRowModule_2_io_H_wire_below_22 ),
       .io_H_wire_below_21( ArrayRowModule_2_io_H_wire_below_21 ),
       .io_H_wire_below_20( ArrayRowModule_2_io_H_wire_below_20 ),
       .io_H_wire_below_19( ArrayRowModule_2_io_H_wire_below_19 ),
       .io_H_wire_below_18( ArrayRowModule_2_io_H_wire_below_18 ),
       .io_H_wire_below_17( ArrayRowModule_2_io_H_wire_below_17 ),
       .io_H_wire_below_16( ArrayRowModule_2_io_H_wire_below_16 ),
       .io_H_wire_below_15( ArrayRowModule_2_io_H_wire_below_15 ),
       .io_H_wire_below_14( ArrayRowModule_2_io_H_wire_below_14 ),
       .io_H_wire_below_13( ArrayRowModule_2_io_H_wire_below_13 ),
       .io_H_wire_below_12( ArrayRowModule_2_io_H_wire_below_12 ),
       .io_H_wire_below_11( ArrayRowModule_2_io_H_wire_below_11 ),
       .io_H_wire_below_10( ArrayRowModule_2_io_H_wire_below_10 ),
       .io_H_wire_below_9( ArrayRowModule_2_io_H_wire_below_9 ),
       .io_H_wire_below_8( ArrayRowModule_2_io_H_wire_below_8 ),
       .io_H_wire_below_7( ArrayRowModule_2_io_H_wire_below_7 ),
       .io_H_wire_below_6( ArrayRowModule_2_io_H_wire_below_6 ),
       .io_H_wire_below_5( ArrayRowModule_2_io_H_wire_below_5 ),
       .io_H_wire_below_4( ArrayRowModule_2_io_H_wire_below_4 ),
       .io_H_wire_below_3( ArrayRowModule_2_io_H_wire_below_3 ),
       .io_H_wire_below_2( ArrayRowModule_2_io_H_wire_below_2 ),
       .io_H_wire_below_1( ArrayRowModule_2_io_H_wire_below_1 ),
       .io_H_wire_below_0( ArrayRowModule_2_io_H_wire_below_0 ),
       .io_row_en( T1473 ),
       //.io_config_or_load(  )
       //.io_D_or_Z(  )
       .io_mem_bus_out_23( ArrayRowModule_2_io_mem_bus_out_23 ),
       .io_mem_bus_out_22( ArrayRowModule_2_io_mem_bus_out_22 ),
       .io_mem_bus_out_21( ArrayRowModule_2_io_mem_bus_out_21 ),
       .io_mem_bus_out_20( ArrayRowModule_2_io_mem_bus_out_20 ),
       .io_mem_bus_out_19( ArrayRowModule_2_io_mem_bus_out_19 ),
       .io_mem_bus_out_18( ArrayRowModule_2_io_mem_bus_out_18 ),
       .io_mem_bus_out_17( ArrayRowModule_2_io_mem_bus_out_17 ),
       .io_mem_bus_out_16( ArrayRowModule_2_io_mem_bus_out_16 ),
       .io_mem_bus_out_15( ArrayRowModule_2_io_mem_bus_out_15 ),
       .io_mem_bus_out_14( ArrayRowModule_2_io_mem_bus_out_14 ),
       .io_mem_bus_out_13( ArrayRowModule_2_io_mem_bus_out_13 ),
       .io_mem_bus_out_12( ArrayRowModule_2_io_mem_bus_out_12 ),
       .io_mem_bus_out_11( ArrayRowModule_2_io_mem_bus_out_11 ),
       .io_mem_bus_out_10( ArrayRowModule_2_io_mem_bus_out_10 ),
       .io_mem_bus_out_9( ArrayRowModule_2_io_mem_bus_out_9 ),
       .io_mem_bus_out_8( ArrayRowModule_2_io_mem_bus_out_8 ),
       .io_mem_bus_out_7( ArrayRowModule_2_io_mem_bus_out_7 ),
       .io_mem_bus_out_6( ArrayRowModule_2_io_mem_bus_out_6 ),
       .io_mem_bus_out_5( ArrayRowModule_2_io_mem_bus_out_5 ),
       .io_mem_bus_out_4( ArrayRowModule_2_io_mem_bus_out_4 ),
       .io_mem_bus_out_3( ArrayRowModule_2_io_mem_bus_out_3 ),
       .io_mem_bus_out_2( ArrayRowModule_2_io_mem_bus_out_2 ),
       .io_mem_bus_out_1( ArrayRowModule_2_io_mem_bus_out_1 ),
       .io_mem_bus_out_0( ArrayRowModule_2_io_mem_bus_out_0 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ArrayRowModule_2.io_config_or_load = {1{$random}};
    assign ArrayRowModule_2.io_D_or_Z = {1{$random}};
    assign ArrayRowModule_2.io_mem_bus_out_23 = {1{$random}};
// synthesis translate_on
`endif
  ArrayRowModule ArrayRowModule_3(.clk(clk), .reset(reset),
       .io_V_wire_in_367( VwireModule_io_VwirePorts_3_22_15_out ),
       .io_V_wire_in_366( VwireModule_io_VwirePorts_3_22_14_out ),
       .io_V_wire_in_365( VwireModule_io_VwirePorts_3_22_13_out ),
       .io_V_wire_in_364( VwireModule_io_VwirePorts_3_22_12_out ),
       .io_V_wire_in_363( VwireModule_io_VwirePorts_3_22_11_out ),
       .io_V_wire_in_362( VwireModule_io_VwirePorts_3_22_10_out ),
       .io_V_wire_in_361( VwireModule_io_VwirePorts_3_22_9_out ),
       .io_V_wire_in_360( VwireModule_io_VwirePorts_3_22_8_out ),
       .io_V_wire_in_359( VwireModule_io_VwirePorts_3_22_7_out ),
       .io_V_wire_in_358( VwireModule_io_VwirePorts_3_22_6_out ),
       .io_V_wire_in_357( VwireModule_io_VwirePorts_3_22_5_out ),
       .io_V_wire_in_356( VwireModule_io_VwirePorts_3_22_4_out ),
       .io_V_wire_in_355( VwireModule_io_VwirePorts_3_22_3_out ),
       .io_V_wire_in_354( VwireModule_io_VwirePorts_3_22_2_out ),
       .io_V_wire_in_353( VwireModule_io_VwirePorts_3_22_1_out ),
       .io_V_wire_in_352( VwireModule_io_VwirePorts_3_22_0_out ),
       .io_V_wire_in_351( VwireModule_io_VwirePorts_3_21_15_out ),
       .io_V_wire_in_350( VwireModule_io_VwirePorts_3_21_14_out ),
       .io_V_wire_in_349( VwireModule_io_VwirePorts_3_21_13_out ),
       .io_V_wire_in_348( VwireModule_io_VwirePorts_3_21_12_out ),
       .io_V_wire_in_347( VwireModule_io_VwirePorts_3_21_11_out ),
       .io_V_wire_in_346( VwireModule_io_VwirePorts_3_21_10_out ),
       .io_V_wire_in_345( VwireModule_io_VwirePorts_3_21_9_out ),
       .io_V_wire_in_344( VwireModule_io_VwirePorts_3_21_8_out ),
       .io_V_wire_in_343( VwireModule_io_VwirePorts_3_21_7_out ),
       .io_V_wire_in_342( VwireModule_io_VwirePorts_3_21_6_out ),
       .io_V_wire_in_341( VwireModule_io_VwirePorts_3_21_5_out ),
       .io_V_wire_in_340( VwireModule_io_VwirePorts_3_21_4_out ),
       .io_V_wire_in_339( VwireModule_io_VwirePorts_3_21_3_out ),
       .io_V_wire_in_338( VwireModule_io_VwirePorts_3_21_2_out ),
       .io_V_wire_in_337( VwireModule_io_VwirePorts_3_21_1_out ),
       .io_V_wire_in_336( VwireModule_io_VwirePorts_3_21_0_out ),
       .io_V_wire_in_335( VwireModule_io_VwirePorts_3_20_15_out ),
       .io_V_wire_in_334( VwireModule_io_VwirePorts_3_20_14_out ),
       .io_V_wire_in_333( VwireModule_io_VwirePorts_3_20_13_out ),
       .io_V_wire_in_332( VwireModule_io_VwirePorts_3_20_12_out ),
       .io_V_wire_in_331( VwireModule_io_VwirePorts_3_20_11_out ),
       .io_V_wire_in_330( VwireModule_io_VwirePorts_3_20_10_out ),
       .io_V_wire_in_329( VwireModule_io_VwirePorts_3_20_9_out ),
       .io_V_wire_in_328( VwireModule_io_VwirePorts_3_20_8_out ),
       .io_V_wire_in_327( VwireModule_io_VwirePorts_3_20_7_out ),
       .io_V_wire_in_326( VwireModule_io_VwirePorts_3_20_6_out ),
       .io_V_wire_in_325( VwireModule_io_VwirePorts_3_20_5_out ),
       .io_V_wire_in_324( VwireModule_io_VwirePorts_3_20_4_out ),
       .io_V_wire_in_323( VwireModule_io_VwirePorts_3_20_3_out ),
       .io_V_wire_in_322( VwireModule_io_VwirePorts_3_20_2_out ),
       .io_V_wire_in_321( VwireModule_io_VwirePorts_3_20_1_out ),
       .io_V_wire_in_320( VwireModule_io_VwirePorts_3_20_0_out ),
       .io_V_wire_in_319( VwireModule_io_VwirePorts_3_19_15_out ),
       .io_V_wire_in_318( VwireModule_io_VwirePorts_3_19_14_out ),
       .io_V_wire_in_317( VwireModule_io_VwirePorts_3_19_13_out ),
       .io_V_wire_in_316( VwireModule_io_VwirePorts_3_19_12_out ),
       .io_V_wire_in_315( VwireModule_io_VwirePorts_3_19_11_out ),
       .io_V_wire_in_314( VwireModule_io_VwirePorts_3_19_10_out ),
       .io_V_wire_in_313( VwireModule_io_VwirePorts_3_19_9_out ),
       .io_V_wire_in_312( VwireModule_io_VwirePorts_3_19_8_out ),
       .io_V_wire_in_311( VwireModule_io_VwirePorts_3_19_7_out ),
       .io_V_wire_in_310( VwireModule_io_VwirePorts_3_19_6_out ),
       .io_V_wire_in_309( VwireModule_io_VwirePorts_3_19_5_out ),
       .io_V_wire_in_308( VwireModule_io_VwirePorts_3_19_4_out ),
       .io_V_wire_in_307( VwireModule_io_VwirePorts_3_19_3_out ),
       .io_V_wire_in_306( VwireModule_io_VwirePorts_3_19_2_out ),
       .io_V_wire_in_305( VwireModule_io_VwirePorts_3_19_1_out ),
       .io_V_wire_in_304( VwireModule_io_VwirePorts_3_19_0_out ),
       .io_V_wire_in_303( VwireModule_io_VwirePorts_3_18_15_out ),
       .io_V_wire_in_302( VwireModule_io_VwirePorts_3_18_14_out ),
       .io_V_wire_in_301( VwireModule_io_VwirePorts_3_18_13_out ),
       .io_V_wire_in_300( VwireModule_io_VwirePorts_3_18_12_out ),
       .io_V_wire_in_299( VwireModule_io_VwirePorts_3_18_11_out ),
       .io_V_wire_in_298( VwireModule_io_VwirePorts_3_18_10_out ),
       .io_V_wire_in_297( VwireModule_io_VwirePorts_3_18_9_out ),
       .io_V_wire_in_296( VwireModule_io_VwirePorts_3_18_8_out ),
       .io_V_wire_in_295( VwireModule_io_VwirePorts_3_18_7_out ),
       .io_V_wire_in_294( VwireModule_io_VwirePorts_3_18_6_out ),
       .io_V_wire_in_293( VwireModule_io_VwirePorts_3_18_5_out ),
       .io_V_wire_in_292( VwireModule_io_VwirePorts_3_18_4_out ),
       .io_V_wire_in_291( VwireModule_io_VwirePorts_3_18_3_out ),
       .io_V_wire_in_290( VwireModule_io_VwirePorts_3_18_2_out ),
       .io_V_wire_in_289( VwireModule_io_VwirePorts_3_18_1_out ),
       .io_V_wire_in_288( VwireModule_io_VwirePorts_3_18_0_out ),
       .io_V_wire_in_287( VwireModule_io_VwirePorts_3_17_15_out ),
       .io_V_wire_in_286( VwireModule_io_VwirePorts_3_17_14_out ),
       .io_V_wire_in_285( VwireModule_io_VwirePorts_3_17_13_out ),
       .io_V_wire_in_284( VwireModule_io_VwirePorts_3_17_12_out ),
       .io_V_wire_in_283( VwireModule_io_VwirePorts_3_17_11_out ),
       .io_V_wire_in_282( VwireModule_io_VwirePorts_3_17_10_out ),
       .io_V_wire_in_281( VwireModule_io_VwirePorts_3_17_9_out ),
       .io_V_wire_in_280( VwireModule_io_VwirePorts_3_17_8_out ),
       .io_V_wire_in_279( VwireModule_io_VwirePorts_3_17_7_out ),
       .io_V_wire_in_278( VwireModule_io_VwirePorts_3_17_6_out ),
       .io_V_wire_in_277( VwireModule_io_VwirePorts_3_17_5_out ),
       .io_V_wire_in_276( VwireModule_io_VwirePorts_3_17_4_out ),
       .io_V_wire_in_275( VwireModule_io_VwirePorts_3_17_3_out ),
       .io_V_wire_in_274( VwireModule_io_VwirePorts_3_17_2_out ),
       .io_V_wire_in_273( VwireModule_io_VwirePorts_3_17_1_out ),
       .io_V_wire_in_272( VwireModule_io_VwirePorts_3_17_0_out ),
       .io_V_wire_in_271( VwireModule_io_VwirePorts_3_16_15_out ),
       .io_V_wire_in_270( VwireModule_io_VwirePorts_3_16_14_out ),
       .io_V_wire_in_269( VwireModule_io_VwirePorts_3_16_13_out ),
       .io_V_wire_in_268( VwireModule_io_VwirePorts_3_16_12_out ),
       .io_V_wire_in_267( VwireModule_io_VwirePorts_3_16_11_out ),
       .io_V_wire_in_266( VwireModule_io_VwirePorts_3_16_10_out ),
       .io_V_wire_in_265( VwireModule_io_VwirePorts_3_16_9_out ),
       .io_V_wire_in_264( VwireModule_io_VwirePorts_3_16_8_out ),
       .io_V_wire_in_263( VwireModule_io_VwirePorts_3_16_7_out ),
       .io_V_wire_in_262( VwireModule_io_VwirePorts_3_16_6_out ),
       .io_V_wire_in_261( VwireModule_io_VwirePorts_3_16_5_out ),
       .io_V_wire_in_260( VwireModule_io_VwirePorts_3_16_4_out ),
       .io_V_wire_in_259( VwireModule_io_VwirePorts_3_16_3_out ),
       .io_V_wire_in_258( VwireModule_io_VwirePorts_3_16_2_out ),
       .io_V_wire_in_257( VwireModule_io_VwirePorts_3_16_1_out ),
       .io_V_wire_in_256( VwireModule_io_VwirePorts_3_16_0_out ),
       .io_V_wire_in_255( VwireModule_io_VwirePorts_3_15_15_out ),
       .io_V_wire_in_254( VwireModule_io_VwirePorts_3_15_14_out ),
       .io_V_wire_in_253( VwireModule_io_VwirePorts_3_15_13_out ),
       .io_V_wire_in_252( VwireModule_io_VwirePorts_3_15_12_out ),
       .io_V_wire_in_251( VwireModule_io_VwirePorts_3_15_11_out ),
       .io_V_wire_in_250( VwireModule_io_VwirePorts_3_15_10_out ),
       .io_V_wire_in_249( VwireModule_io_VwirePorts_3_15_9_out ),
       .io_V_wire_in_248( VwireModule_io_VwirePorts_3_15_8_out ),
       .io_V_wire_in_247( VwireModule_io_VwirePorts_3_15_7_out ),
       .io_V_wire_in_246( VwireModule_io_VwirePorts_3_15_6_out ),
       .io_V_wire_in_245( VwireModule_io_VwirePorts_3_15_5_out ),
       .io_V_wire_in_244( VwireModule_io_VwirePorts_3_15_4_out ),
       .io_V_wire_in_243( VwireModule_io_VwirePorts_3_15_3_out ),
       .io_V_wire_in_242( VwireModule_io_VwirePorts_3_15_2_out ),
       .io_V_wire_in_241( VwireModule_io_VwirePorts_3_15_1_out ),
       .io_V_wire_in_240( VwireModule_io_VwirePorts_3_15_0_out ),
       .io_V_wire_in_239( VwireModule_io_VwirePorts_3_14_15_out ),
       .io_V_wire_in_238( VwireModule_io_VwirePorts_3_14_14_out ),
       .io_V_wire_in_237( VwireModule_io_VwirePorts_3_14_13_out ),
       .io_V_wire_in_236( VwireModule_io_VwirePorts_3_14_12_out ),
       .io_V_wire_in_235( VwireModule_io_VwirePorts_3_14_11_out ),
       .io_V_wire_in_234( VwireModule_io_VwirePorts_3_14_10_out ),
       .io_V_wire_in_233( VwireModule_io_VwirePorts_3_14_9_out ),
       .io_V_wire_in_232( VwireModule_io_VwirePorts_3_14_8_out ),
       .io_V_wire_in_231( VwireModule_io_VwirePorts_3_14_7_out ),
       .io_V_wire_in_230( VwireModule_io_VwirePorts_3_14_6_out ),
       .io_V_wire_in_229( VwireModule_io_VwirePorts_3_14_5_out ),
       .io_V_wire_in_228( VwireModule_io_VwirePorts_3_14_4_out ),
       .io_V_wire_in_227( VwireModule_io_VwirePorts_3_14_3_out ),
       .io_V_wire_in_226( VwireModule_io_VwirePorts_3_14_2_out ),
       .io_V_wire_in_225( VwireModule_io_VwirePorts_3_14_1_out ),
       .io_V_wire_in_224( VwireModule_io_VwirePorts_3_14_0_out ),
       .io_V_wire_in_223( VwireModule_io_VwirePorts_3_13_15_out ),
       .io_V_wire_in_222( VwireModule_io_VwirePorts_3_13_14_out ),
       .io_V_wire_in_221( VwireModule_io_VwirePorts_3_13_13_out ),
       .io_V_wire_in_220( VwireModule_io_VwirePorts_3_13_12_out ),
       .io_V_wire_in_219( VwireModule_io_VwirePorts_3_13_11_out ),
       .io_V_wire_in_218( VwireModule_io_VwirePorts_3_13_10_out ),
       .io_V_wire_in_217( VwireModule_io_VwirePorts_3_13_9_out ),
       .io_V_wire_in_216( VwireModule_io_VwirePorts_3_13_8_out ),
       .io_V_wire_in_215( VwireModule_io_VwirePorts_3_13_7_out ),
       .io_V_wire_in_214( VwireModule_io_VwirePorts_3_13_6_out ),
       .io_V_wire_in_213( VwireModule_io_VwirePorts_3_13_5_out ),
       .io_V_wire_in_212( VwireModule_io_VwirePorts_3_13_4_out ),
       .io_V_wire_in_211( VwireModule_io_VwirePorts_3_13_3_out ),
       .io_V_wire_in_210( VwireModule_io_VwirePorts_3_13_2_out ),
       .io_V_wire_in_209( VwireModule_io_VwirePorts_3_13_1_out ),
       .io_V_wire_in_208( VwireModule_io_VwirePorts_3_13_0_out ),
       .io_V_wire_in_207( VwireModule_io_VwirePorts_3_12_15_out ),
       .io_V_wire_in_206( VwireModule_io_VwirePorts_3_12_14_out ),
       .io_V_wire_in_205( VwireModule_io_VwirePorts_3_12_13_out ),
       .io_V_wire_in_204( VwireModule_io_VwirePorts_3_12_12_out ),
       .io_V_wire_in_203( VwireModule_io_VwirePorts_3_12_11_out ),
       .io_V_wire_in_202( VwireModule_io_VwirePorts_3_12_10_out ),
       .io_V_wire_in_201( VwireModule_io_VwirePorts_3_12_9_out ),
       .io_V_wire_in_200( VwireModule_io_VwirePorts_3_12_8_out ),
       .io_V_wire_in_199( VwireModule_io_VwirePorts_3_12_7_out ),
       .io_V_wire_in_198( VwireModule_io_VwirePorts_3_12_6_out ),
       .io_V_wire_in_197( VwireModule_io_VwirePorts_3_12_5_out ),
       .io_V_wire_in_196( VwireModule_io_VwirePorts_3_12_4_out ),
       .io_V_wire_in_195( VwireModule_io_VwirePorts_3_12_3_out ),
       .io_V_wire_in_194( VwireModule_io_VwirePorts_3_12_2_out ),
       .io_V_wire_in_193( VwireModule_io_VwirePorts_3_12_1_out ),
       .io_V_wire_in_192( VwireModule_io_VwirePorts_3_12_0_out ),
       .io_V_wire_in_191( VwireModule_io_VwirePorts_3_11_15_out ),
       .io_V_wire_in_190( VwireModule_io_VwirePorts_3_11_14_out ),
       .io_V_wire_in_189( VwireModule_io_VwirePorts_3_11_13_out ),
       .io_V_wire_in_188( VwireModule_io_VwirePorts_3_11_12_out ),
       .io_V_wire_in_187( VwireModule_io_VwirePorts_3_11_11_out ),
       .io_V_wire_in_186( VwireModule_io_VwirePorts_3_11_10_out ),
       .io_V_wire_in_185( VwireModule_io_VwirePorts_3_11_9_out ),
       .io_V_wire_in_184( VwireModule_io_VwirePorts_3_11_8_out ),
       .io_V_wire_in_183( VwireModule_io_VwirePorts_3_11_7_out ),
       .io_V_wire_in_182( VwireModule_io_VwirePorts_3_11_6_out ),
       .io_V_wire_in_181( VwireModule_io_VwirePorts_3_11_5_out ),
       .io_V_wire_in_180( VwireModule_io_VwirePorts_3_11_4_out ),
       .io_V_wire_in_179( VwireModule_io_VwirePorts_3_11_3_out ),
       .io_V_wire_in_178( VwireModule_io_VwirePorts_3_11_2_out ),
       .io_V_wire_in_177( VwireModule_io_VwirePorts_3_11_1_out ),
       .io_V_wire_in_176( VwireModule_io_VwirePorts_3_11_0_out ),
       .io_V_wire_in_175( VwireModule_io_VwirePorts_3_10_15_out ),
       .io_V_wire_in_174( VwireModule_io_VwirePorts_3_10_14_out ),
       .io_V_wire_in_173( VwireModule_io_VwirePorts_3_10_13_out ),
       .io_V_wire_in_172( VwireModule_io_VwirePorts_3_10_12_out ),
       .io_V_wire_in_171( VwireModule_io_VwirePorts_3_10_11_out ),
       .io_V_wire_in_170( VwireModule_io_VwirePorts_3_10_10_out ),
       .io_V_wire_in_169( VwireModule_io_VwirePorts_3_10_9_out ),
       .io_V_wire_in_168( VwireModule_io_VwirePorts_3_10_8_out ),
       .io_V_wire_in_167( VwireModule_io_VwirePorts_3_10_7_out ),
       .io_V_wire_in_166( VwireModule_io_VwirePorts_3_10_6_out ),
       .io_V_wire_in_165( VwireModule_io_VwirePorts_3_10_5_out ),
       .io_V_wire_in_164( VwireModule_io_VwirePorts_3_10_4_out ),
       .io_V_wire_in_163( VwireModule_io_VwirePorts_3_10_3_out ),
       .io_V_wire_in_162( VwireModule_io_VwirePorts_3_10_2_out ),
       .io_V_wire_in_161( VwireModule_io_VwirePorts_3_10_1_out ),
       .io_V_wire_in_160( VwireModule_io_VwirePorts_3_10_0_out ),
       .io_V_wire_in_159( VwireModule_io_VwirePorts_3_9_15_out ),
       .io_V_wire_in_158( VwireModule_io_VwirePorts_3_9_14_out ),
       .io_V_wire_in_157( VwireModule_io_VwirePorts_3_9_13_out ),
       .io_V_wire_in_156( VwireModule_io_VwirePorts_3_9_12_out ),
       .io_V_wire_in_155( VwireModule_io_VwirePorts_3_9_11_out ),
       .io_V_wire_in_154( VwireModule_io_VwirePorts_3_9_10_out ),
       .io_V_wire_in_153( VwireModule_io_VwirePorts_3_9_9_out ),
       .io_V_wire_in_152( VwireModule_io_VwirePorts_3_9_8_out ),
       .io_V_wire_in_151( VwireModule_io_VwirePorts_3_9_7_out ),
       .io_V_wire_in_150( VwireModule_io_VwirePorts_3_9_6_out ),
       .io_V_wire_in_149( VwireModule_io_VwirePorts_3_9_5_out ),
       .io_V_wire_in_148( VwireModule_io_VwirePorts_3_9_4_out ),
       .io_V_wire_in_147( VwireModule_io_VwirePorts_3_9_3_out ),
       .io_V_wire_in_146( VwireModule_io_VwirePorts_3_9_2_out ),
       .io_V_wire_in_145( VwireModule_io_VwirePorts_3_9_1_out ),
       .io_V_wire_in_144( VwireModule_io_VwirePorts_3_9_0_out ),
       .io_V_wire_in_143( VwireModule_io_VwirePorts_3_8_15_out ),
       .io_V_wire_in_142( VwireModule_io_VwirePorts_3_8_14_out ),
       .io_V_wire_in_141( VwireModule_io_VwirePorts_3_8_13_out ),
       .io_V_wire_in_140( VwireModule_io_VwirePorts_3_8_12_out ),
       .io_V_wire_in_139( VwireModule_io_VwirePorts_3_8_11_out ),
       .io_V_wire_in_138( VwireModule_io_VwirePorts_3_8_10_out ),
       .io_V_wire_in_137( VwireModule_io_VwirePorts_3_8_9_out ),
       .io_V_wire_in_136( VwireModule_io_VwirePorts_3_8_8_out ),
       .io_V_wire_in_135( VwireModule_io_VwirePorts_3_8_7_out ),
       .io_V_wire_in_134( VwireModule_io_VwirePorts_3_8_6_out ),
       .io_V_wire_in_133( VwireModule_io_VwirePorts_3_8_5_out ),
       .io_V_wire_in_132( VwireModule_io_VwirePorts_3_8_4_out ),
       .io_V_wire_in_131( VwireModule_io_VwirePorts_3_8_3_out ),
       .io_V_wire_in_130( VwireModule_io_VwirePorts_3_8_2_out ),
       .io_V_wire_in_129( VwireModule_io_VwirePorts_3_8_1_out ),
       .io_V_wire_in_128( VwireModule_io_VwirePorts_3_8_0_out ),
       .io_V_wire_in_127( VwireModule_io_VwirePorts_3_7_15_out ),
       .io_V_wire_in_126( VwireModule_io_VwirePorts_3_7_14_out ),
       .io_V_wire_in_125( VwireModule_io_VwirePorts_3_7_13_out ),
       .io_V_wire_in_124( VwireModule_io_VwirePorts_3_7_12_out ),
       .io_V_wire_in_123( VwireModule_io_VwirePorts_3_7_11_out ),
       .io_V_wire_in_122( VwireModule_io_VwirePorts_3_7_10_out ),
       .io_V_wire_in_121( VwireModule_io_VwirePorts_3_7_9_out ),
       .io_V_wire_in_120( VwireModule_io_VwirePorts_3_7_8_out ),
       .io_V_wire_in_119( VwireModule_io_VwirePorts_3_7_7_out ),
       .io_V_wire_in_118( VwireModule_io_VwirePorts_3_7_6_out ),
       .io_V_wire_in_117( VwireModule_io_VwirePorts_3_7_5_out ),
       .io_V_wire_in_116( VwireModule_io_VwirePorts_3_7_4_out ),
       .io_V_wire_in_115( VwireModule_io_VwirePorts_3_7_3_out ),
       .io_V_wire_in_114( VwireModule_io_VwirePorts_3_7_2_out ),
       .io_V_wire_in_113( VwireModule_io_VwirePorts_3_7_1_out ),
       .io_V_wire_in_112( VwireModule_io_VwirePorts_3_7_0_out ),
       .io_V_wire_in_111( VwireModule_io_VwirePorts_3_6_15_out ),
       .io_V_wire_in_110( VwireModule_io_VwirePorts_3_6_14_out ),
       .io_V_wire_in_109( VwireModule_io_VwirePorts_3_6_13_out ),
       .io_V_wire_in_108( VwireModule_io_VwirePorts_3_6_12_out ),
       .io_V_wire_in_107( VwireModule_io_VwirePorts_3_6_11_out ),
       .io_V_wire_in_106( VwireModule_io_VwirePorts_3_6_10_out ),
       .io_V_wire_in_105( VwireModule_io_VwirePorts_3_6_9_out ),
       .io_V_wire_in_104( VwireModule_io_VwirePorts_3_6_8_out ),
       .io_V_wire_in_103( VwireModule_io_VwirePorts_3_6_7_out ),
       .io_V_wire_in_102( VwireModule_io_VwirePorts_3_6_6_out ),
       .io_V_wire_in_101( VwireModule_io_VwirePorts_3_6_5_out ),
       .io_V_wire_in_100( VwireModule_io_VwirePorts_3_6_4_out ),
       .io_V_wire_in_99( VwireModule_io_VwirePorts_3_6_3_out ),
       .io_V_wire_in_98( VwireModule_io_VwirePorts_3_6_2_out ),
       .io_V_wire_in_97( VwireModule_io_VwirePorts_3_6_1_out ),
       .io_V_wire_in_96( VwireModule_io_VwirePorts_3_6_0_out ),
       .io_V_wire_in_95( VwireModule_io_VwirePorts_3_5_15_out ),
       .io_V_wire_in_94( VwireModule_io_VwirePorts_3_5_14_out ),
       .io_V_wire_in_93( VwireModule_io_VwirePorts_3_5_13_out ),
       .io_V_wire_in_92( VwireModule_io_VwirePorts_3_5_12_out ),
       .io_V_wire_in_91( VwireModule_io_VwirePorts_3_5_11_out ),
       .io_V_wire_in_90( VwireModule_io_VwirePorts_3_5_10_out ),
       .io_V_wire_in_89( VwireModule_io_VwirePorts_3_5_9_out ),
       .io_V_wire_in_88( VwireModule_io_VwirePorts_3_5_8_out ),
       .io_V_wire_in_87( VwireModule_io_VwirePorts_3_5_7_out ),
       .io_V_wire_in_86( VwireModule_io_VwirePorts_3_5_6_out ),
       .io_V_wire_in_85( VwireModule_io_VwirePorts_3_5_5_out ),
       .io_V_wire_in_84( VwireModule_io_VwirePorts_3_5_4_out ),
       .io_V_wire_in_83( VwireModule_io_VwirePorts_3_5_3_out ),
       .io_V_wire_in_82( VwireModule_io_VwirePorts_3_5_2_out ),
       .io_V_wire_in_81( VwireModule_io_VwirePorts_3_5_1_out ),
       .io_V_wire_in_80( VwireModule_io_VwirePorts_3_5_0_out ),
       .io_V_wire_in_79( VwireModule_io_VwirePorts_3_4_15_out ),
       .io_V_wire_in_78( VwireModule_io_VwirePorts_3_4_14_out ),
       .io_V_wire_in_77( VwireModule_io_VwirePorts_3_4_13_out ),
       .io_V_wire_in_76( VwireModule_io_VwirePorts_3_4_12_out ),
       .io_V_wire_in_75( VwireModule_io_VwirePorts_3_4_11_out ),
       .io_V_wire_in_74( VwireModule_io_VwirePorts_3_4_10_out ),
       .io_V_wire_in_73( VwireModule_io_VwirePorts_3_4_9_out ),
       .io_V_wire_in_72( VwireModule_io_VwirePorts_3_4_8_out ),
       .io_V_wire_in_71( VwireModule_io_VwirePorts_3_4_7_out ),
       .io_V_wire_in_70( VwireModule_io_VwirePorts_3_4_6_out ),
       .io_V_wire_in_69( VwireModule_io_VwirePorts_3_4_5_out ),
       .io_V_wire_in_68( VwireModule_io_VwirePorts_3_4_4_out ),
       .io_V_wire_in_67( VwireModule_io_VwirePorts_3_4_3_out ),
       .io_V_wire_in_66( VwireModule_io_VwirePorts_3_4_2_out ),
       .io_V_wire_in_65( VwireModule_io_VwirePorts_3_4_1_out ),
       .io_V_wire_in_64( VwireModule_io_VwirePorts_3_4_0_out ),
       .io_V_wire_in_63( VwireModule_io_VwirePorts_3_3_15_out ),
       .io_V_wire_in_62( VwireModule_io_VwirePorts_3_3_14_out ),
       .io_V_wire_in_61( VwireModule_io_VwirePorts_3_3_13_out ),
       .io_V_wire_in_60( VwireModule_io_VwirePorts_3_3_12_out ),
       .io_V_wire_in_59( VwireModule_io_VwirePorts_3_3_11_out ),
       .io_V_wire_in_58( VwireModule_io_VwirePorts_3_3_10_out ),
       .io_V_wire_in_57( VwireModule_io_VwirePorts_3_3_9_out ),
       .io_V_wire_in_56( VwireModule_io_VwirePorts_3_3_8_out ),
       .io_V_wire_in_55( VwireModule_io_VwirePorts_3_3_7_out ),
       .io_V_wire_in_54( VwireModule_io_VwirePorts_3_3_6_out ),
       .io_V_wire_in_53( VwireModule_io_VwirePorts_3_3_5_out ),
       .io_V_wire_in_52( VwireModule_io_VwirePorts_3_3_4_out ),
       .io_V_wire_in_51( VwireModule_io_VwirePorts_3_3_3_out ),
       .io_V_wire_in_50( VwireModule_io_VwirePorts_3_3_2_out ),
       .io_V_wire_in_49( VwireModule_io_VwirePorts_3_3_1_out ),
       .io_V_wire_in_48( VwireModule_io_VwirePorts_3_3_0_out ),
       .io_V_wire_in_47( VwireModule_io_VwirePorts_3_2_15_out ),
       .io_V_wire_in_46( VwireModule_io_VwirePorts_3_2_14_out ),
       .io_V_wire_in_45( VwireModule_io_VwirePorts_3_2_13_out ),
       .io_V_wire_in_44( VwireModule_io_VwirePorts_3_2_12_out ),
       .io_V_wire_in_43( VwireModule_io_VwirePorts_3_2_11_out ),
       .io_V_wire_in_42( VwireModule_io_VwirePorts_3_2_10_out ),
       .io_V_wire_in_41( VwireModule_io_VwirePorts_3_2_9_out ),
       .io_V_wire_in_40( VwireModule_io_VwirePorts_3_2_8_out ),
       .io_V_wire_in_39( VwireModule_io_VwirePorts_3_2_7_out ),
       .io_V_wire_in_38( VwireModule_io_VwirePorts_3_2_6_out ),
       .io_V_wire_in_37( VwireModule_io_VwirePorts_3_2_5_out ),
       .io_V_wire_in_36( VwireModule_io_VwirePorts_3_2_4_out ),
       .io_V_wire_in_35( VwireModule_io_VwirePorts_3_2_3_out ),
       .io_V_wire_in_34( VwireModule_io_VwirePorts_3_2_2_out ),
       .io_V_wire_in_33( VwireModule_io_VwirePorts_3_2_1_out ),
       .io_V_wire_in_32( VwireModule_io_VwirePorts_3_2_0_out ),
       .io_V_wire_in_31( VwireModule_io_VwirePorts_3_1_15_out ),
       .io_V_wire_in_30( VwireModule_io_VwirePorts_3_1_14_out ),
       .io_V_wire_in_29( VwireModule_io_VwirePorts_3_1_13_out ),
       .io_V_wire_in_28( VwireModule_io_VwirePorts_3_1_12_out ),
       .io_V_wire_in_27( VwireModule_io_VwirePorts_3_1_11_out ),
       .io_V_wire_in_26( VwireModule_io_VwirePorts_3_1_10_out ),
       .io_V_wire_in_25( VwireModule_io_VwirePorts_3_1_9_out ),
       .io_V_wire_in_24( VwireModule_io_VwirePorts_3_1_8_out ),
       .io_V_wire_in_23( VwireModule_io_VwirePorts_3_1_7_out ),
       .io_V_wire_in_22( VwireModule_io_VwirePorts_3_1_6_out ),
       .io_V_wire_in_21( VwireModule_io_VwirePorts_3_1_5_out ),
       .io_V_wire_in_20( VwireModule_io_VwirePorts_3_1_4_out ),
       .io_V_wire_in_19( VwireModule_io_VwirePorts_3_1_3_out ),
       .io_V_wire_in_18( VwireModule_io_VwirePorts_3_1_2_out ),
       .io_V_wire_in_17( VwireModule_io_VwirePorts_3_1_1_out ),
       .io_V_wire_in_16( VwireModule_io_VwirePorts_3_1_0_out ),
       .io_V_wire_in_15( VwireModule_io_VwirePorts_3_0_15_out ),
       .io_V_wire_in_14( VwireModule_io_VwirePorts_3_0_14_out ),
       .io_V_wire_in_13( VwireModule_io_VwirePorts_3_0_13_out ),
       .io_V_wire_in_12( VwireModule_io_VwirePorts_3_0_12_out ),
       .io_V_wire_in_11( VwireModule_io_VwirePorts_3_0_11_out ),
       .io_V_wire_in_10( VwireModule_io_VwirePorts_3_0_10_out ),
       .io_V_wire_in_9( VwireModule_io_VwirePorts_3_0_9_out ),
       .io_V_wire_in_8( VwireModule_io_VwirePorts_3_0_8_out ),
       .io_V_wire_in_7( VwireModule_io_VwirePorts_3_0_7_out ),
       .io_V_wire_in_6( VwireModule_io_VwirePorts_3_0_6_out ),
       .io_V_wire_in_5( VwireModule_io_VwirePorts_3_0_5_out ),
       .io_V_wire_in_4( VwireModule_io_VwirePorts_3_0_4_out ),
       .io_V_wire_in_3( VwireModule_io_VwirePorts_3_0_3_out ),
       .io_V_wire_in_2( VwireModule_io_VwirePorts_3_0_2_out ),
       .io_V_wire_in_1( VwireModule_io_VwirePorts_3_0_1_out ),
       .io_V_wire_in_0( VwireModule_io_VwirePorts_3_0_0_out ),
       .io_V_wire_out_367( ArrayRowModule_3_io_V_wire_out_367 ),
       .io_V_wire_out_366( ArrayRowModule_3_io_V_wire_out_366 ),
       .io_V_wire_out_365( ArrayRowModule_3_io_V_wire_out_365 ),
       .io_V_wire_out_364( ArrayRowModule_3_io_V_wire_out_364 ),
       .io_V_wire_out_363( ArrayRowModule_3_io_V_wire_out_363 ),
       .io_V_wire_out_362( ArrayRowModule_3_io_V_wire_out_362 ),
       .io_V_wire_out_361( ArrayRowModule_3_io_V_wire_out_361 ),
       .io_V_wire_out_360( ArrayRowModule_3_io_V_wire_out_360 ),
       .io_V_wire_out_359( ArrayRowModule_3_io_V_wire_out_359 ),
       .io_V_wire_out_358( ArrayRowModule_3_io_V_wire_out_358 ),
       .io_V_wire_out_357( ArrayRowModule_3_io_V_wire_out_357 ),
       .io_V_wire_out_356( ArrayRowModule_3_io_V_wire_out_356 ),
       .io_V_wire_out_355( ArrayRowModule_3_io_V_wire_out_355 ),
       .io_V_wire_out_354( ArrayRowModule_3_io_V_wire_out_354 ),
       .io_V_wire_out_353( ArrayRowModule_3_io_V_wire_out_353 ),
       .io_V_wire_out_352( ArrayRowModule_3_io_V_wire_out_352 ),
       .io_V_wire_out_351( ArrayRowModule_3_io_V_wire_out_351 ),
       .io_V_wire_out_350( ArrayRowModule_3_io_V_wire_out_350 ),
       .io_V_wire_out_349( ArrayRowModule_3_io_V_wire_out_349 ),
       .io_V_wire_out_348( ArrayRowModule_3_io_V_wire_out_348 ),
       .io_V_wire_out_347( ArrayRowModule_3_io_V_wire_out_347 ),
       .io_V_wire_out_346( ArrayRowModule_3_io_V_wire_out_346 ),
       .io_V_wire_out_345( ArrayRowModule_3_io_V_wire_out_345 ),
       .io_V_wire_out_344( ArrayRowModule_3_io_V_wire_out_344 ),
       .io_V_wire_out_343( ArrayRowModule_3_io_V_wire_out_343 ),
       .io_V_wire_out_342( ArrayRowModule_3_io_V_wire_out_342 ),
       .io_V_wire_out_341( ArrayRowModule_3_io_V_wire_out_341 ),
       .io_V_wire_out_340( ArrayRowModule_3_io_V_wire_out_340 ),
       .io_V_wire_out_339( ArrayRowModule_3_io_V_wire_out_339 ),
       .io_V_wire_out_338( ArrayRowModule_3_io_V_wire_out_338 ),
       .io_V_wire_out_337( ArrayRowModule_3_io_V_wire_out_337 ),
       .io_V_wire_out_336( ArrayRowModule_3_io_V_wire_out_336 ),
       .io_V_wire_out_335( ArrayRowModule_3_io_V_wire_out_335 ),
       .io_V_wire_out_334( ArrayRowModule_3_io_V_wire_out_334 ),
       .io_V_wire_out_333( ArrayRowModule_3_io_V_wire_out_333 ),
       .io_V_wire_out_332( ArrayRowModule_3_io_V_wire_out_332 ),
       .io_V_wire_out_331( ArrayRowModule_3_io_V_wire_out_331 ),
       .io_V_wire_out_330( ArrayRowModule_3_io_V_wire_out_330 ),
       .io_V_wire_out_329( ArrayRowModule_3_io_V_wire_out_329 ),
       .io_V_wire_out_328( ArrayRowModule_3_io_V_wire_out_328 ),
       .io_V_wire_out_327( ArrayRowModule_3_io_V_wire_out_327 ),
       .io_V_wire_out_326( ArrayRowModule_3_io_V_wire_out_326 ),
       .io_V_wire_out_325( ArrayRowModule_3_io_V_wire_out_325 ),
       .io_V_wire_out_324( ArrayRowModule_3_io_V_wire_out_324 ),
       .io_V_wire_out_323( ArrayRowModule_3_io_V_wire_out_323 ),
       .io_V_wire_out_322( ArrayRowModule_3_io_V_wire_out_322 ),
       .io_V_wire_out_321( ArrayRowModule_3_io_V_wire_out_321 ),
       .io_V_wire_out_320( ArrayRowModule_3_io_V_wire_out_320 ),
       .io_V_wire_out_319( ArrayRowModule_3_io_V_wire_out_319 ),
       .io_V_wire_out_318( ArrayRowModule_3_io_V_wire_out_318 ),
       .io_V_wire_out_317( ArrayRowModule_3_io_V_wire_out_317 ),
       .io_V_wire_out_316( ArrayRowModule_3_io_V_wire_out_316 ),
       .io_V_wire_out_315( ArrayRowModule_3_io_V_wire_out_315 ),
       .io_V_wire_out_314( ArrayRowModule_3_io_V_wire_out_314 ),
       .io_V_wire_out_313( ArrayRowModule_3_io_V_wire_out_313 ),
       .io_V_wire_out_312( ArrayRowModule_3_io_V_wire_out_312 ),
       .io_V_wire_out_311( ArrayRowModule_3_io_V_wire_out_311 ),
       .io_V_wire_out_310( ArrayRowModule_3_io_V_wire_out_310 ),
       .io_V_wire_out_309( ArrayRowModule_3_io_V_wire_out_309 ),
       .io_V_wire_out_308( ArrayRowModule_3_io_V_wire_out_308 ),
       .io_V_wire_out_307( ArrayRowModule_3_io_V_wire_out_307 ),
       .io_V_wire_out_306( ArrayRowModule_3_io_V_wire_out_306 ),
       .io_V_wire_out_305( ArrayRowModule_3_io_V_wire_out_305 ),
       .io_V_wire_out_304( ArrayRowModule_3_io_V_wire_out_304 ),
       .io_V_wire_out_303( ArrayRowModule_3_io_V_wire_out_303 ),
       .io_V_wire_out_302( ArrayRowModule_3_io_V_wire_out_302 ),
       .io_V_wire_out_301( ArrayRowModule_3_io_V_wire_out_301 ),
       .io_V_wire_out_300( ArrayRowModule_3_io_V_wire_out_300 ),
       .io_V_wire_out_299( ArrayRowModule_3_io_V_wire_out_299 ),
       .io_V_wire_out_298( ArrayRowModule_3_io_V_wire_out_298 ),
       .io_V_wire_out_297( ArrayRowModule_3_io_V_wire_out_297 ),
       .io_V_wire_out_296( ArrayRowModule_3_io_V_wire_out_296 ),
       .io_V_wire_out_295( ArrayRowModule_3_io_V_wire_out_295 ),
       .io_V_wire_out_294( ArrayRowModule_3_io_V_wire_out_294 ),
       .io_V_wire_out_293( ArrayRowModule_3_io_V_wire_out_293 ),
       .io_V_wire_out_292( ArrayRowModule_3_io_V_wire_out_292 ),
       .io_V_wire_out_291( ArrayRowModule_3_io_V_wire_out_291 ),
       .io_V_wire_out_290( ArrayRowModule_3_io_V_wire_out_290 ),
       .io_V_wire_out_289( ArrayRowModule_3_io_V_wire_out_289 ),
       .io_V_wire_out_288( ArrayRowModule_3_io_V_wire_out_288 ),
       .io_V_wire_out_287( ArrayRowModule_3_io_V_wire_out_287 ),
       .io_V_wire_out_286( ArrayRowModule_3_io_V_wire_out_286 ),
       .io_V_wire_out_285( ArrayRowModule_3_io_V_wire_out_285 ),
       .io_V_wire_out_284( ArrayRowModule_3_io_V_wire_out_284 ),
       .io_V_wire_out_283( ArrayRowModule_3_io_V_wire_out_283 ),
       .io_V_wire_out_282( ArrayRowModule_3_io_V_wire_out_282 ),
       .io_V_wire_out_281( ArrayRowModule_3_io_V_wire_out_281 ),
       .io_V_wire_out_280( ArrayRowModule_3_io_V_wire_out_280 ),
       .io_V_wire_out_279( ArrayRowModule_3_io_V_wire_out_279 ),
       .io_V_wire_out_278( ArrayRowModule_3_io_V_wire_out_278 ),
       .io_V_wire_out_277( ArrayRowModule_3_io_V_wire_out_277 ),
       .io_V_wire_out_276( ArrayRowModule_3_io_V_wire_out_276 ),
       .io_V_wire_out_275( ArrayRowModule_3_io_V_wire_out_275 ),
       .io_V_wire_out_274( ArrayRowModule_3_io_V_wire_out_274 ),
       .io_V_wire_out_273( ArrayRowModule_3_io_V_wire_out_273 ),
       .io_V_wire_out_272( ArrayRowModule_3_io_V_wire_out_272 ),
       .io_V_wire_out_271( ArrayRowModule_3_io_V_wire_out_271 ),
       .io_V_wire_out_270( ArrayRowModule_3_io_V_wire_out_270 ),
       .io_V_wire_out_269( ArrayRowModule_3_io_V_wire_out_269 ),
       .io_V_wire_out_268( ArrayRowModule_3_io_V_wire_out_268 ),
       .io_V_wire_out_267( ArrayRowModule_3_io_V_wire_out_267 ),
       .io_V_wire_out_266( ArrayRowModule_3_io_V_wire_out_266 ),
       .io_V_wire_out_265( ArrayRowModule_3_io_V_wire_out_265 ),
       .io_V_wire_out_264( ArrayRowModule_3_io_V_wire_out_264 ),
       .io_V_wire_out_263( ArrayRowModule_3_io_V_wire_out_263 ),
       .io_V_wire_out_262( ArrayRowModule_3_io_V_wire_out_262 ),
       .io_V_wire_out_261( ArrayRowModule_3_io_V_wire_out_261 ),
       .io_V_wire_out_260( ArrayRowModule_3_io_V_wire_out_260 ),
       .io_V_wire_out_259( ArrayRowModule_3_io_V_wire_out_259 ),
       .io_V_wire_out_258( ArrayRowModule_3_io_V_wire_out_258 ),
       .io_V_wire_out_257( ArrayRowModule_3_io_V_wire_out_257 ),
       .io_V_wire_out_256( ArrayRowModule_3_io_V_wire_out_256 ),
       .io_V_wire_out_255( ArrayRowModule_3_io_V_wire_out_255 ),
       .io_V_wire_out_254( ArrayRowModule_3_io_V_wire_out_254 ),
       .io_V_wire_out_253( ArrayRowModule_3_io_V_wire_out_253 ),
       .io_V_wire_out_252( ArrayRowModule_3_io_V_wire_out_252 ),
       .io_V_wire_out_251( ArrayRowModule_3_io_V_wire_out_251 ),
       .io_V_wire_out_250( ArrayRowModule_3_io_V_wire_out_250 ),
       .io_V_wire_out_249( ArrayRowModule_3_io_V_wire_out_249 ),
       .io_V_wire_out_248( ArrayRowModule_3_io_V_wire_out_248 ),
       .io_V_wire_out_247( ArrayRowModule_3_io_V_wire_out_247 ),
       .io_V_wire_out_246( ArrayRowModule_3_io_V_wire_out_246 ),
       .io_V_wire_out_245( ArrayRowModule_3_io_V_wire_out_245 ),
       .io_V_wire_out_244( ArrayRowModule_3_io_V_wire_out_244 ),
       .io_V_wire_out_243( ArrayRowModule_3_io_V_wire_out_243 ),
       .io_V_wire_out_242( ArrayRowModule_3_io_V_wire_out_242 ),
       .io_V_wire_out_241( ArrayRowModule_3_io_V_wire_out_241 ),
       .io_V_wire_out_240( ArrayRowModule_3_io_V_wire_out_240 ),
       .io_V_wire_out_239( ArrayRowModule_3_io_V_wire_out_239 ),
       .io_V_wire_out_238( ArrayRowModule_3_io_V_wire_out_238 ),
       .io_V_wire_out_237( ArrayRowModule_3_io_V_wire_out_237 ),
       .io_V_wire_out_236( ArrayRowModule_3_io_V_wire_out_236 ),
       .io_V_wire_out_235( ArrayRowModule_3_io_V_wire_out_235 ),
       .io_V_wire_out_234( ArrayRowModule_3_io_V_wire_out_234 ),
       .io_V_wire_out_233( ArrayRowModule_3_io_V_wire_out_233 ),
       .io_V_wire_out_232( ArrayRowModule_3_io_V_wire_out_232 ),
       .io_V_wire_out_231( ArrayRowModule_3_io_V_wire_out_231 ),
       .io_V_wire_out_230( ArrayRowModule_3_io_V_wire_out_230 ),
       .io_V_wire_out_229( ArrayRowModule_3_io_V_wire_out_229 ),
       .io_V_wire_out_228( ArrayRowModule_3_io_V_wire_out_228 ),
       .io_V_wire_out_227( ArrayRowModule_3_io_V_wire_out_227 ),
       .io_V_wire_out_226( ArrayRowModule_3_io_V_wire_out_226 ),
       .io_V_wire_out_225( ArrayRowModule_3_io_V_wire_out_225 ),
       .io_V_wire_out_224( ArrayRowModule_3_io_V_wire_out_224 ),
       .io_V_wire_out_223( ArrayRowModule_3_io_V_wire_out_223 ),
       .io_V_wire_out_222( ArrayRowModule_3_io_V_wire_out_222 ),
       .io_V_wire_out_221( ArrayRowModule_3_io_V_wire_out_221 ),
       .io_V_wire_out_220( ArrayRowModule_3_io_V_wire_out_220 ),
       .io_V_wire_out_219( ArrayRowModule_3_io_V_wire_out_219 ),
       .io_V_wire_out_218( ArrayRowModule_3_io_V_wire_out_218 ),
       .io_V_wire_out_217( ArrayRowModule_3_io_V_wire_out_217 ),
       .io_V_wire_out_216( ArrayRowModule_3_io_V_wire_out_216 ),
       .io_V_wire_out_215( ArrayRowModule_3_io_V_wire_out_215 ),
       .io_V_wire_out_214( ArrayRowModule_3_io_V_wire_out_214 ),
       .io_V_wire_out_213( ArrayRowModule_3_io_V_wire_out_213 ),
       .io_V_wire_out_212( ArrayRowModule_3_io_V_wire_out_212 ),
       .io_V_wire_out_211( ArrayRowModule_3_io_V_wire_out_211 ),
       .io_V_wire_out_210( ArrayRowModule_3_io_V_wire_out_210 ),
       .io_V_wire_out_209( ArrayRowModule_3_io_V_wire_out_209 ),
       .io_V_wire_out_208( ArrayRowModule_3_io_V_wire_out_208 ),
       .io_V_wire_out_207( ArrayRowModule_3_io_V_wire_out_207 ),
       .io_V_wire_out_206( ArrayRowModule_3_io_V_wire_out_206 ),
       .io_V_wire_out_205( ArrayRowModule_3_io_V_wire_out_205 ),
       .io_V_wire_out_204( ArrayRowModule_3_io_V_wire_out_204 ),
       .io_V_wire_out_203( ArrayRowModule_3_io_V_wire_out_203 ),
       .io_V_wire_out_202( ArrayRowModule_3_io_V_wire_out_202 ),
       .io_V_wire_out_201( ArrayRowModule_3_io_V_wire_out_201 ),
       .io_V_wire_out_200( ArrayRowModule_3_io_V_wire_out_200 ),
       .io_V_wire_out_199( ArrayRowModule_3_io_V_wire_out_199 ),
       .io_V_wire_out_198( ArrayRowModule_3_io_V_wire_out_198 ),
       .io_V_wire_out_197( ArrayRowModule_3_io_V_wire_out_197 ),
       .io_V_wire_out_196( ArrayRowModule_3_io_V_wire_out_196 ),
       .io_V_wire_out_195( ArrayRowModule_3_io_V_wire_out_195 ),
       .io_V_wire_out_194( ArrayRowModule_3_io_V_wire_out_194 ),
       .io_V_wire_out_193( ArrayRowModule_3_io_V_wire_out_193 ),
       .io_V_wire_out_192( ArrayRowModule_3_io_V_wire_out_192 ),
       .io_V_wire_out_191( ArrayRowModule_3_io_V_wire_out_191 ),
       .io_V_wire_out_190( ArrayRowModule_3_io_V_wire_out_190 ),
       .io_V_wire_out_189( ArrayRowModule_3_io_V_wire_out_189 ),
       .io_V_wire_out_188( ArrayRowModule_3_io_V_wire_out_188 ),
       .io_V_wire_out_187( ArrayRowModule_3_io_V_wire_out_187 ),
       .io_V_wire_out_186( ArrayRowModule_3_io_V_wire_out_186 ),
       .io_V_wire_out_185( ArrayRowModule_3_io_V_wire_out_185 ),
       .io_V_wire_out_184( ArrayRowModule_3_io_V_wire_out_184 ),
       .io_V_wire_out_183( ArrayRowModule_3_io_V_wire_out_183 ),
       .io_V_wire_out_182( ArrayRowModule_3_io_V_wire_out_182 ),
       .io_V_wire_out_181( ArrayRowModule_3_io_V_wire_out_181 ),
       .io_V_wire_out_180( ArrayRowModule_3_io_V_wire_out_180 ),
       .io_V_wire_out_179( ArrayRowModule_3_io_V_wire_out_179 ),
       .io_V_wire_out_178( ArrayRowModule_3_io_V_wire_out_178 ),
       .io_V_wire_out_177( ArrayRowModule_3_io_V_wire_out_177 ),
       .io_V_wire_out_176( ArrayRowModule_3_io_V_wire_out_176 ),
       .io_V_wire_out_175( ArrayRowModule_3_io_V_wire_out_175 ),
       .io_V_wire_out_174( ArrayRowModule_3_io_V_wire_out_174 ),
       .io_V_wire_out_173( ArrayRowModule_3_io_V_wire_out_173 ),
       .io_V_wire_out_172( ArrayRowModule_3_io_V_wire_out_172 ),
       .io_V_wire_out_171( ArrayRowModule_3_io_V_wire_out_171 ),
       .io_V_wire_out_170( ArrayRowModule_3_io_V_wire_out_170 ),
       .io_V_wire_out_169( ArrayRowModule_3_io_V_wire_out_169 ),
       .io_V_wire_out_168( ArrayRowModule_3_io_V_wire_out_168 ),
       .io_V_wire_out_167( ArrayRowModule_3_io_V_wire_out_167 ),
       .io_V_wire_out_166( ArrayRowModule_3_io_V_wire_out_166 ),
       .io_V_wire_out_165( ArrayRowModule_3_io_V_wire_out_165 ),
       .io_V_wire_out_164( ArrayRowModule_3_io_V_wire_out_164 ),
       .io_V_wire_out_163( ArrayRowModule_3_io_V_wire_out_163 ),
       .io_V_wire_out_162( ArrayRowModule_3_io_V_wire_out_162 ),
       .io_V_wire_out_161( ArrayRowModule_3_io_V_wire_out_161 ),
       .io_V_wire_out_160( ArrayRowModule_3_io_V_wire_out_160 ),
       .io_V_wire_out_159( ArrayRowModule_3_io_V_wire_out_159 ),
       .io_V_wire_out_158( ArrayRowModule_3_io_V_wire_out_158 ),
       .io_V_wire_out_157( ArrayRowModule_3_io_V_wire_out_157 ),
       .io_V_wire_out_156( ArrayRowModule_3_io_V_wire_out_156 ),
       .io_V_wire_out_155( ArrayRowModule_3_io_V_wire_out_155 ),
       .io_V_wire_out_154( ArrayRowModule_3_io_V_wire_out_154 ),
       .io_V_wire_out_153( ArrayRowModule_3_io_V_wire_out_153 ),
       .io_V_wire_out_152( ArrayRowModule_3_io_V_wire_out_152 ),
       .io_V_wire_out_151( ArrayRowModule_3_io_V_wire_out_151 ),
       .io_V_wire_out_150( ArrayRowModule_3_io_V_wire_out_150 ),
       .io_V_wire_out_149( ArrayRowModule_3_io_V_wire_out_149 ),
       .io_V_wire_out_148( ArrayRowModule_3_io_V_wire_out_148 ),
       .io_V_wire_out_147( ArrayRowModule_3_io_V_wire_out_147 ),
       .io_V_wire_out_146( ArrayRowModule_3_io_V_wire_out_146 ),
       .io_V_wire_out_145( ArrayRowModule_3_io_V_wire_out_145 ),
       .io_V_wire_out_144( ArrayRowModule_3_io_V_wire_out_144 ),
       .io_V_wire_out_143( ArrayRowModule_3_io_V_wire_out_143 ),
       .io_V_wire_out_142( ArrayRowModule_3_io_V_wire_out_142 ),
       .io_V_wire_out_141( ArrayRowModule_3_io_V_wire_out_141 ),
       .io_V_wire_out_140( ArrayRowModule_3_io_V_wire_out_140 ),
       .io_V_wire_out_139( ArrayRowModule_3_io_V_wire_out_139 ),
       .io_V_wire_out_138( ArrayRowModule_3_io_V_wire_out_138 ),
       .io_V_wire_out_137( ArrayRowModule_3_io_V_wire_out_137 ),
       .io_V_wire_out_136( ArrayRowModule_3_io_V_wire_out_136 ),
       .io_V_wire_out_135( ArrayRowModule_3_io_V_wire_out_135 ),
       .io_V_wire_out_134( ArrayRowModule_3_io_V_wire_out_134 ),
       .io_V_wire_out_133( ArrayRowModule_3_io_V_wire_out_133 ),
       .io_V_wire_out_132( ArrayRowModule_3_io_V_wire_out_132 ),
       .io_V_wire_out_131( ArrayRowModule_3_io_V_wire_out_131 ),
       .io_V_wire_out_130( ArrayRowModule_3_io_V_wire_out_130 ),
       .io_V_wire_out_129( ArrayRowModule_3_io_V_wire_out_129 ),
       .io_V_wire_out_128( ArrayRowModule_3_io_V_wire_out_128 ),
       .io_V_wire_out_127( ArrayRowModule_3_io_V_wire_out_127 ),
       .io_V_wire_out_126( ArrayRowModule_3_io_V_wire_out_126 ),
       .io_V_wire_out_125( ArrayRowModule_3_io_V_wire_out_125 ),
       .io_V_wire_out_124( ArrayRowModule_3_io_V_wire_out_124 ),
       .io_V_wire_out_123( ArrayRowModule_3_io_V_wire_out_123 ),
       .io_V_wire_out_122( ArrayRowModule_3_io_V_wire_out_122 ),
       .io_V_wire_out_121( ArrayRowModule_3_io_V_wire_out_121 ),
       .io_V_wire_out_120( ArrayRowModule_3_io_V_wire_out_120 ),
       .io_V_wire_out_119( ArrayRowModule_3_io_V_wire_out_119 ),
       .io_V_wire_out_118( ArrayRowModule_3_io_V_wire_out_118 ),
       .io_V_wire_out_117( ArrayRowModule_3_io_V_wire_out_117 ),
       .io_V_wire_out_116( ArrayRowModule_3_io_V_wire_out_116 ),
       .io_V_wire_out_115( ArrayRowModule_3_io_V_wire_out_115 ),
       .io_V_wire_out_114( ArrayRowModule_3_io_V_wire_out_114 ),
       .io_V_wire_out_113( ArrayRowModule_3_io_V_wire_out_113 ),
       .io_V_wire_out_112( ArrayRowModule_3_io_V_wire_out_112 ),
       .io_V_wire_out_111( ArrayRowModule_3_io_V_wire_out_111 ),
       .io_V_wire_out_110( ArrayRowModule_3_io_V_wire_out_110 ),
       .io_V_wire_out_109( ArrayRowModule_3_io_V_wire_out_109 ),
       .io_V_wire_out_108( ArrayRowModule_3_io_V_wire_out_108 ),
       .io_V_wire_out_107( ArrayRowModule_3_io_V_wire_out_107 ),
       .io_V_wire_out_106( ArrayRowModule_3_io_V_wire_out_106 ),
       .io_V_wire_out_105( ArrayRowModule_3_io_V_wire_out_105 ),
       .io_V_wire_out_104( ArrayRowModule_3_io_V_wire_out_104 ),
       .io_V_wire_out_103( ArrayRowModule_3_io_V_wire_out_103 ),
       .io_V_wire_out_102( ArrayRowModule_3_io_V_wire_out_102 ),
       .io_V_wire_out_101( ArrayRowModule_3_io_V_wire_out_101 ),
       .io_V_wire_out_100( ArrayRowModule_3_io_V_wire_out_100 ),
       .io_V_wire_out_99( ArrayRowModule_3_io_V_wire_out_99 ),
       .io_V_wire_out_98( ArrayRowModule_3_io_V_wire_out_98 ),
       .io_V_wire_out_97( ArrayRowModule_3_io_V_wire_out_97 ),
       .io_V_wire_out_96( ArrayRowModule_3_io_V_wire_out_96 ),
       .io_V_wire_out_95( ArrayRowModule_3_io_V_wire_out_95 ),
       .io_V_wire_out_94( ArrayRowModule_3_io_V_wire_out_94 ),
       .io_V_wire_out_93( ArrayRowModule_3_io_V_wire_out_93 ),
       .io_V_wire_out_92( ArrayRowModule_3_io_V_wire_out_92 ),
       .io_V_wire_out_91( ArrayRowModule_3_io_V_wire_out_91 ),
       .io_V_wire_out_90( ArrayRowModule_3_io_V_wire_out_90 ),
       .io_V_wire_out_89( ArrayRowModule_3_io_V_wire_out_89 ),
       .io_V_wire_out_88( ArrayRowModule_3_io_V_wire_out_88 ),
       .io_V_wire_out_87( ArrayRowModule_3_io_V_wire_out_87 ),
       .io_V_wire_out_86( ArrayRowModule_3_io_V_wire_out_86 ),
       .io_V_wire_out_85( ArrayRowModule_3_io_V_wire_out_85 ),
       .io_V_wire_out_84( ArrayRowModule_3_io_V_wire_out_84 ),
       .io_V_wire_out_83( ArrayRowModule_3_io_V_wire_out_83 ),
       .io_V_wire_out_82( ArrayRowModule_3_io_V_wire_out_82 ),
       .io_V_wire_out_81( ArrayRowModule_3_io_V_wire_out_81 ),
       .io_V_wire_out_80( ArrayRowModule_3_io_V_wire_out_80 ),
       .io_V_wire_out_79( ArrayRowModule_3_io_V_wire_out_79 ),
       .io_V_wire_out_78( ArrayRowModule_3_io_V_wire_out_78 ),
       .io_V_wire_out_77( ArrayRowModule_3_io_V_wire_out_77 ),
       .io_V_wire_out_76( ArrayRowModule_3_io_V_wire_out_76 ),
       .io_V_wire_out_75( ArrayRowModule_3_io_V_wire_out_75 ),
       .io_V_wire_out_74( ArrayRowModule_3_io_V_wire_out_74 ),
       .io_V_wire_out_73( ArrayRowModule_3_io_V_wire_out_73 ),
       .io_V_wire_out_72( ArrayRowModule_3_io_V_wire_out_72 ),
       .io_V_wire_out_71( ArrayRowModule_3_io_V_wire_out_71 ),
       .io_V_wire_out_70( ArrayRowModule_3_io_V_wire_out_70 ),
       .io_V_wire_out_69( ArrayRowModule_3_io_V_wire_out_69 ),
       .io_V_wire_out_68( ArrayRowModule_3_io_V_wire_out_68 ),
       .io_V_wire_out_67( ArrayRowModule_3_io_V_wire_out_67 ),
       .io_V_wire_out_66( ArrayRowModule_3_io_V_wire_out_66 ),
       .io_V_wire_out_65( ArrayRowModule_3_io_V_wire_out_65 ),
       .io_V_wire_out_64( ArrayRowModule_3_io_V_wire_out_64 ),
       .io_V_wire_out_63( ArrayRowModule_3_io_V_wire_out_63 ),
       .io_V_wire_out_62( ArrayRowModule_3_io_V_wire_out_62 ),
       .io_V_wire_out_61( ArrayRowModule_3_io_V_wire_out_61 ),
       .io_V_wire_out_60( ArrayRowModule_3_io_V_wire_out_60 ),
       .io_V_wire_out_59( ArrayRowModule_3_io_V_wire_out_59 ),
       .io_V_wire_out_58( ArrayRowModule_3_io_V_wire_out_58 ),
       .io_V_wire_out_57( ArrayRowModule_3_io_V_wire_out_57 ),
       .io_V_wire_out_56( ArrayRowModule_3_io_V_wire_out_56 ),
       .io_V_wire_out_55( ArrayRowModule_3_io_V_wire_out_55 ),
       .io_V_wire_out_54( ArrayRowModule_3_io_V_wire_out_54 ),
       .io_V_wire_out_53( ArrayRowModule_3_io_V_wire_out_53 ),
       .io_V_wire_out_52( ArrayRowModule_3_io_V_wire_out_52 ),
       .io_V_wire_out_51( ArrayRowModule_3_io_V_wire_out_51 ),
       .io_V_wire_out_50( ArrayRowModule_3_io_V_wire_out_50 ),
       .io_V_wire_out_49( ArrayRowModule_3_io_V_wire_out_49 ),
       .io_V_wire_out_48( ArrayRowModule_3_io_V_wire_out_48 ),
       .io_V_wire_out_47( ArrayRowModule_3_io_V_wire_out_47 ),
       .io_V_wire_out_46( ArrayRowModule_3_io_V_wire_out_46 ),
       .io_V_wire_out_45( ArrayRowModule_3_io_V_wire_out_45 ),
       .io_V_wire_out_44( ArrayRowModule_3_io_V_wire_out_44 ),
       .io_V_wire_out_43( ArrayRowModule_3_io_V_wire_out_43 ),
       .io_V_wire_out_42( ArrayRowModule_3_io_V_wire_out_42 ),
       .io_V_wire_out_41( ArrayRowModule_3_io_V_wire_out_41 ),
       .io_V_wire_out_40( ArrayRowModule_3_io_V_wire_out_40 ),
       .io_V_wire_out_39( ArrayRowModule_3_io_V_wire_out_39 ),
       .io_V_wire_out_38( ArrayRowModule_3_io_V_wire_out_38 ),
       .io_V_wire_out_37( ArrayRowModule_3_io_V_wire_out_37 ),
       .io_V_wire_out_36( ArrayRowModule_3_io_V_wire_out_36 ),
       .io_V_wire_out_35( ArrayRowModule_3_io_V_wire_out_35 ),
       .io_V_wire_out_34( ArrayRowModule_3_io_V_wire_out_34 ),
       .io_V_wire_out_33( ArrayRowModule_3_io_V_wire_out_33 ),
       .io_V_wire_out_32( ArrayRowModule_3_io_V_wire_out_32 ),
       .io_V_wire_out_31( ArrayRowModule_3_io_V_wire_out_31 ),
       .io_V_wire_out_30( ArrayRowModule_3_io_V_wire_out_30 ),
       .io_V_wire_out_29( ArrayRowModule_3_io_V_wire_out_29 ),
       .io_V_wire_out_28( ArrayRowModule_3_io_V_wire_out_28 ),
       .io_V_wire_out_27( ArrayRowModule_3_io_V_wire_out_27 ),
       .io_V_wire_out_26( ArrayRowModule_3_io_V_wire_out_26 ),
       .io_V_wire_out_25( ArrayRowModule_3_io_V_wire_out_25 ),
       .io_V_wire_out_24( ArrayRowModule_3_io_V_wire_out_24 ),
       .io_V_wire_out_23( ArrayRowModule_3_io_V_wire_out_23 ),
       .io_V_wire_out_22( ArrayRowModule_3_io_V_wire_out_22 ),
       .io_V_wire_out_21( ArrayRowModule_3_io_V_wire_out_21 ),
       .io_V_wire_out_20( ArrayRowModule_3_io_V_wire_out_20 ),
       .io_V_wire_out_19( ArrayRowModule_3_io_V_wire_out_19 ),
       .io_V_wire_out_18( ArrayRowModule_3_io_V_wire_out_18 ),
       .io_V_wire_out_17( ArrayRowModule_3_io_V_wire_out_17 ),
       .io_V_wire_out_16( ArrayRowModule_3_io_V_wire_out_16 ),
       .io_V_wire_out_15( ArrayRowModule_3_io_V_wire_out_15 ),
       .io_V_wire_out_14( ArrayRowModule_3_io_V_wire_out_14 ),
       .io_V_wire_out_13( ArrayRowModule_3_io_V_wire_out_13 ),
       .io_V_wire_out_12( ArrayRowModule_3_io_V_wire_out_12 ),
       .io_V_wire_out_11( ArrayRowModule_3_io_V_wire_out_11 ),
       .io_V_wire_out_10( ArrayRowModule_3_io_V_wire_out_10 ),
       .io_V_wire_out_9( ArrayRowModule_3_io_V_wire_out_9 ),
       .io_V_wire_out_8( ArrayRowModule_3_io_V_wire_out_8 ),
       .io_V_wire_out_7( ArrayRowModule_3_io_V_wire_out_7 ),
       .io_V_wire_out_6( ArrayRowModule_3_io_V_wire_out_6 ),
       .io_V_wire_out_5( ArrayRowModule_3_io_V_wire_out_5 ),
       .io_V_wire_out_4( ArrayRowModule_3_io_V_wire_out_4 ),
       .io_V_wire_out_3( ArrayRowModule_3_io_V_wire_out_3 ),
       .io_V_wire_out_2( ArrayRowModule_3_io_V_wire_out_2 ),
       .io_V_wire_out_1( ArrayRowModule_3_io_V_wire_out_1 ),
       .io_V_wire_out_0( ArrayRowModule_3_io_V_wire_out_0 ),
       .io_V_wire_en_22( ArrayRowModule_3_io_V_wire_en_22 ),
       .io_V_wire_en_21( ArrayRowModule_3_io_V_wire_en_21 ),
       .io_V_wire_en_20( ArrayRowModule_3_io_V_wire_en_20 ),
       .io_V_wire_en_19( ArrayRowModule_3_io_V_wire_en_19 ),
       .io_V_wire_en_18( ArrayRowModule_3_io_V_wire_en_18 ),
       .io_V_wire_en_17( ArrayRowModule_3_io_V_wire_en_17 ),
       .io_V_wire_en_16( ArrayRowModule_3_io_V_wire_en_16 ),
       .io_V_wire_en_15( ArrayRowModule_3_io_V_wire_en_15 ),
       .io_V_wire_en_14( ArrayRowModule_3_io_V_wire_en_14 ),
       .io_V_wire_en_13( ArrayRowModule_3_io_V_wire_en_13 ),
       .io_V_wire_en_12( ArrayRowModule_3_io_V_wire_en_12 ),
       .io_V_wire_en_11( ArrayRowModule_3_io_V_wire_en_11 ),
       .io_V_wire_en_10( ArrayRowModule_3_io_V_wire_en_10 ),
       .io_V_wire_en_9( ArrayRowModule_3_io_V_wire_en_9 ),
       .io_V_wire_en_8( ArrayRowModule_3_io_V_wire_en_8 ),
       .io_V_wire_en_7( ArrayRowModule_3_io_V_wire_en_7 ),
       .io_V_wire_en_6( ArrayRowModule_3_io_V_wire_en_6 ),
       .io_V_wire_en_5( ArrayRowModule_3_io_V_wire_en_5 ),
       .io_V_wire_en_4( ArrayRowModule_3_io_V_wire_en_4 ),
       .io_V_wire_en_3( ArrayRowModule_3_io_V_wire_en_3 ),
       .io_V_wire_en_2( ArrayRowModule_3_io_V_wire_en_2 ),
       .io_V_wire_en_1( ArrayRowModule_3_io_V_wire_en_1 ),
       .io_V_wire_en_0( ArrayRowModule_3_io_V_wire_en_0 ),
       .io_G_wire_above_3( ArrayRowModule_2_io_G_wire_below_3 ),
       .io_G_wire_above_2( ArrayRowModule_2_io_G_wire_below_2 ),
       .io_G_wire_above_1( ArrayRowModule_2_io_G_wire_below_1 ),
       .io_G_wire_above_0( ArrayRowModule_2_io_G_wire_below_0 ),
       .io_H_wire_above_32( ArrayRowModule_2_io_H_wire_below_32 ),
       .io_H_wire_above_31( ArrayRowModule_2_io_H_wire_below_31 ),
       .io_H_wire_above_30( ArrayRowModule_2_io_H_wire_below_30 ),
       .io_H_wire_above_29( ArrayRowModule_2_io_H_wire_below_29 ),
       .io_H_wire_above_28( ArrayRowModule_2_io_H_wire_below_28 ),
       .io_H_wire_above_27( ArrayRowModule_2_io_H_wire_below_27 ),
       .io_H_wire_above_26( ArrayRowModule_2_io_H_wire_below_26 ),
       .io_H_wire_above_25( ArrayRowModule_2_io_H_wire_below_25 ),
       .io_H_wire_above_24( ArrayRowModule_2_io_H_wire_below_24 ),
       .io_H_wire_above_23( ArrayRowModule_2_io_H_wire_below_23 ),
       .io_H_wire_above_22( ArrayRowModule_2_io_H_wire_below_22 ),
       .io_H_wire_above_21( ArrayRowModule_2_io_H_wire_below_21 ),
       .io_H_wire_above_20( ArrayRowModule_2_io_H_wire_below_20 ),
       .io_H_wire_above_19( ArrayRowModule_2_io_H_wire_below_19 ),
       .io_H_wire_above_18( ArrayRowModule_2_io_H_wire_below_18 ),
       .io_H_wire_above_17( ArrayRowModule_2_io_H_wire_below_17 ),
       .io_H_wire_above_16( ArrayRowModule_2_io_H_wire_below_16 ),
       .io_H_wire_above_15( ArrayRowModule_2_io_H_wire_below_15 ),
       .io_H_wire_above_14( ArrayRowModule_2_io_H_wire_below_14 ),
       .io_H_wire_above_13( ArrayRowModule_2_io_H_wire_below_13 ),
       .io_H_wire_above_12( ArrayRowModule_2_io_H_wire_below_12 ),
       .io_H_wire_above_11( ArrayRowModule_2_io_H_wire_below_11 ),
       .io_H_wire_above_10( ArrayRowModule_2_io_H_wire_below_10 ),
       .io_H_wire_above_9( ArrayRowModule_2_io_H_wire_below_9 ),
       .io_H_wire_above_8( ArrayRowModule_2_io_H_wire_below_8 ),
       .io_H_wire_above_7( ArrayRowModule_2_io_H_wire_below_7 ),
       .io_H_wire_above_6( ArrayRowModule_2_io_H_wire_below_6 ),
       .io_H_wire_above_5( ArrayRowModule_2_io_H_wire_below_5 ),
       .io_H_wire_above_4( ArrayRowModule_2_io_H_wire_below_4 ),
       .io_H_wire_above_3( ArrayRowModule_2_io_H_wire_below_3 ),
       .io_H_wire_above_2( ArrayRowModule_2_io_H_wire_below_2 ),
       .io_H_wire_above_1( ArrayRowModule_2_io_H_wire_below_1 ),
       .io_H_wire_above_0( ArrayRowModule_2_io_H_wire_below_0 ),
       .io_mem_bus_in_23( ArrayRowModule_2_io_mem_bus_out_23 ),
       .io_mem_bus_in_22( ArrayRowModule_2_io_mem_bus_out_22 ),
       .io_mem_bus_in_21( ArrayRowModule_2_io_mem_bus_out_21 ),
       .io_mem_bus_in_20( ArrayRowModule_2_io_mem_bus_out_20 ),
       .io_mem_bus_in_19( ArrayRowModule_2_io_mem_bus_out_19 ),
       .io_mem_bus_in_18( ArrayRowModule_2_io_mem_bus_out_18 ),
       .io_mem_bus_in_17( ArrayRowModule_2_io_mem_bus_out_17 ),
       .io_mem_bus_in_16( ArrayRowModule_2_io_mem_bus_out_16 ),
       .io_mem_bus_in_15( ArrayRowModule_2_io_mem_bus_out_15 ),
       .io_mem_bus_in_14( ArrayRowModule_2_io_mem_bus_out_14 ),
       .io_mem_bus_in_13( ArrayRowModule_2_io_mem_bus_out_13 ),
       .io_mem_bus_in_12( ArrayRowModule_2_io_mem_bus_out_12 ),
       .io_mem_bus_in_11( ArrayRowModule_2_io_mem_bus_out_11 ),
       .io_mem_bus_in_10( ArrayRowModule_2_io_mem_bus_out_10 ),
       .io_mem_bus_in_9( ArrayRowModule_2_io_mem_bus_out_9 ),
       .io_mem_bus_in_8( ArrayRowModule_2_io_mem_bus_out_8 ),
       .io_mem_bus_in_7( ArrayRowModule_2_io_mem_bus_out_7 ),
       .io_mem_bus_in_6( ArrayRowModule_2_io_mem_bus_out_6 ),
       .io_mem_bus_in_5( ArrayRowModule_2_io_mem_bus_out_5 ),
       .io_mem_bus_in_4( ArrayRowModule_2_io_mem_bus_out_4 ),
       .io_mem_bus_in_3( ArrayRowModule_2_io_mem_bus_out_3 ),
       .io_mem_bus_in_2( ArrayRowModule_2_io_mem_bus_out_2 ),
       .io_mem_bus_in_1( ArrayRowModule_2_io_mem_bus_out_1 ),
       .io_mem_bus_in_0( ArrayRowModule_2_io_mem_bus_out_0 ),
       .io_H_out_above_22( ArrayRowModule_2_io_H_out_22 ),
       .io_H_out_above_21( ArrayRowModule_2_io_H_out_21 ),
       .io_H_out_above_20( ArrayRowModule_2_io_H_out_20 ),
       .io_H_out_above_19( ArrayRowModule_2_io_H_out_19 ),
       .io_H_out_above_18( ArrayRowModule_2_io_H_out_18 ),
       .io_H_out_above_17( ArrayRowModule_2_io_H_out_17 ),
       .io_H_out_above_16( ArrayRowModule_2_io_H_out_16 ),
       .io_H_out_above_15( ArrayRowModule_2_io_H_out_15 ),
       .io_H_out_above_14( ArrayRowModule_2_io_H_out_14 ),
       .io_H_out_above_13( ArrayRowModule_2_io_H_out_13 ),
       .io_H_out_above_12( ArrayRowModule_2_io_H_out_12 ),
       .io_H_out_above_11( ArrayRowModule_2_io_H_out_11 ),
       .io_H_out_above_10( ArrayRowModule_2_io_H_out_10 ),
       .io_H_out_above_9( ArrayRowModule_2_io_H_out_9 ),
       .io_H_out_above_8( ArrayRowModule_2_io_H_out_8 ),
       .io_H_out_above_7( ArrayRowModule_2_io_H_out_7 ),
       .io_H_out_above_6( ArrayRowModule_2_io_H_out_6 ),
       .io_H_out_above_5( ArrayRowModule_2_io_H_out_5 ),
       .io_H_out_above_4( ArrayRowModule_2_io_H_out_4 ),
       .io_H_out_above_3( ArrayRowModule_2_io_H_out_3 ),
       .io_H_out_above_2( ArrayRowModule_2_io_H_out_2 ),
       .io_H_out_above_1( ArrayRowModule_2_io_H_out_1 ),
       .io_H_out_above_0( ArrayRowModule_2_io_H_out_0 ),
       //.io_H_out_22(  )
       //.io_H_out_21(  )
       //.io_H_out_20(  )
       //.io_H_out_19(  )
       //.io_H_out_18(  )
       //.io_H_out_17(  )
       //.io_H_out_16(  )
       //.io_H_out_15(  )
       //.io_H_out_14(  )
       //.io_H_out_13(  )
       //.io_H_out_12(  )
       //.io_H_out_11(  )
       //.io_H_out_10(  )
       //.io_H_out_9(  )
       //.io_H_out_8(  )
       //.io_H_out_7(  )
       //.io_H_out_6(  )
       //.io_H_out_5(  )
       //.io_H_out_4(  )
       //.io_H_out_3(  )
       //.io_H_out_2(  )
       //.io_H_out_1(  )
       //.io_H_out_0(  )
       //.io_G_wire_below_3(  )
       //.io_G_wire_below_2(  )
       //.io_G_wire_below_1(  )
       //.io_G_wire_below_0(  )
       //.io_H_wire_below_32(  )
       //.io_H_wire_below_31(  )
       //.io_H_wire_below_30(  )
       //.io_H_wire_below_29(  )
       //.io_H_wire_below_28(  )
       //.io_H_wire_below_27(  )
       //.io_H_wire_below_26(  )
       //.io_H_wire_below_25(  )
       //.io_H_wire_below_24(  )
       //.io_H_wire_below_23(  )
       //.io_H_wire_below_22(  )
       //.io_H_wire_below_21(  )
       //.io_H_wire_below_20(  )
       //.io_H_wire_below_19(  )
       //.io_H_wire_below_18(  )
       //.io_H_wire_below_17(  )
       //.io_H_wire_below_16(  )
       //.io_H_wire_below_15(  )
       //.io_H_wire_below_14(  )
       //.io_H_wire_below_13(  )
       //.io_H_wire_below_12(  )
       //.io_H_wire_below_11(  )
       //.io_H_wire_below_10(  )
       //.io_H_wire_below_9(  )
       //.io_H_wire_below_8(  )
       //.io_H_wire_below_7(  )
       //.io_H_wire_below_6(  )
       //.io_H_wire_below_5(  )
       //.io_H_wire_below_4(  )
       //.io_H_wire_below_3(  )
       //.io_H_wire_below_2(  )
       //.io_H_wire_below_1(  )
       //.io_H_wire_below_0(  )
       .io_row_en( T1472 ),
       //.io_config_or_load(  )
       //.io_D_or_Z(  )
       .io_mem_bus_out_23( ArrayRowModule_3_io_mem_bus_out_23 ),
       .io_mem_bus_out_22( ArrayRowModule_3_io_mem_bus_out_22 ),
       .io_mem_bus_out_21( ArrayRowModule_3_io_mem_bus_out_21 ),
       .io_mem_bus_out_20( ArrayRowModule_3_io_mem_bus_out_20 ),
       .io_mem_bus_out_19( ArrayRowModule_3_io_mem_bus_out_19 ),
       .io_mem_bus_out_18( ArrayRowModule_3_io_mem_bus_out_18 ),
       .io_mem_bus_out_17( ArrayRowModule_3_io_mem_bus_out_17 ),
       .io_mem_bus_out_16( ArrayRowModule_3_io_mem_bus_out_16 ),
       .io_mem_bus_out_15( ArrayRowModule_3_io_mem_bus_out_15 ),
       .io_mem_bus_out_14( ArrayRowModule_3_io_mem_bus_out_14 ),
       .io_mem_bus_out_13( ArrayRowModule_3_io_mem_bus_out_13 ),
       .io_mem_bus_out_12( ArrayRowModule_3_io_mem_bus_out_12 ),
       .io_mem_bus_out_11( ArrayRowModule_3_io_mem_bus_out_11 ),
       .io_mem_bus_out_10( ArrayRowModule_3_io_mem_bus_out_10 ),
       .io_mem_bus_out_9( ArrayRowModule_3_io_mem_bus_out_9 ),
       .io_mem_bus_out_8( ArrayRowModule_3_io_mem_bus_out_8 ),
       .io_mem_bus_out_7( ArrayRowModule_3_io_mem_bus_out_7 ),
       .io_mem_bus_out_6( ArrayRowModule_3_io_mem_bus_out_6 ),
       .io_mem_bus_out_5( ArrayRowModule_3_io_mem_bus_out_5 ),
       .io_mem_bus_out_4( ArrayRowModule_3_io_mem_bus_out_4 ),
       .io_mem_bus_out_3( ArrayRowModule_3_io_mem_bus_out_3 ),
       .io_mem_bus_out_2( ArrayRowModule_3_io_mem_bus_out_2 ),
       .io_mem_bus_out_1( ArrayRowModule_3_io_mem_bus_out_1 ),
       .io_mem_bus_out_0( ArrayRowModule_3_io_mem_bus_out_0 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ArrayRowModule_3.io_config_or_load = {1{$random}};
    assign ArrayRowModule_3.io_D_or_Z = {1{$random}};
    assign ArrayRowModule_3.io_mem_bus_out_23 = {1{$random}};
// synthesis translate_on
`endif
  VwireModule VwireModule(
       .io_VwirePorts_3_22_15_in( ArrayRowModule_3_io_V_wire_out_367 ),
       .io_VwirePorts_3_22_15_en( T1471 ),
       .io_VwirePorts_3_22_15_out( VwireModule_io_VwirePorts_3_22_15_out ),
       .io_VwirePorts_3_22_14_in( ArrayRowModule_3_io_V_wire_out_366 ),
       .io_VwirePorts_3_22_14_en( T1470 ),
       .io_VwirePorts_3_22_14_out( VwireModule_io_VwirePorts_3_22_14_out ),
       .io_VwirePorts_3_22_13_in( ArrayRowModule_3_io_V_wire_out_365 ),
       .io_VwirePorts_3_22_13_en( T1469 ),
       .io_VwirePorts_3_22_13_out( VwireModule_io_VwirePorts_3_22_13_out ),
       .io_VwirePorts_3_22_12_in( ArrayRowModule_3_io_V_wire_out_364 ),
       .io_VwirePorts_3_22_12_en( T1468 ),
       .io_VwirePorts_3_22_12_out( VwireModule_io_VwirePorts_3_22_12_out ),
       .io_VwirePorts_3_22_11_in( ArrayRowModule_3_io_V_wire_out_363 ),
       .io_VwirePorts_3_22_11_en( T1467 ),
       .io_VwirePorts_3_22_11_out( VwireModule_io_VwirePorts_3_22_11_out ),
       .io_VwirePorts_3_22_10_in( ArrayRowModule_3_io_V_wire_out_362 ),
       .io_VwirePorts_3_22_10_en( T1466 ),
       .io_VwirePorts_3_22_10_out( VwireModule_io_VwirePorts_3_22_10_out ),
       .io_VwirePorts_3_22_9_in( ArrayRowModule_3_io_V_wire_out_361 ),
       .io_VwirePorts_3_22_9_en( T1465 ),
       .io_VwirePorts_3_22_9_out( VwireModule_io_VwirePorts_3_22_9_out ),
       .io_VwirePorts_3_22_8_in( ArrayRowModule_3_io_V_wire_out_360 ),
       .io_VwirePorts_3_22_8_en( T1464 ),
       .io_VwirePorts_3_22_8_out( VwireModule_io_VwirePorts_3_22_8_out ),
       .io_VwirePorts_3_22_7_in( ArrayRowModule_3_io_V_wire_out_359 ),
       .io_VwirePorts_3_22_7_en( T1463 ),
       .io_VwirePorts_3_22_7_out( VwireModule_io_VwirePorts_3_22_7_out ),
       .io_VwirePorts_3_22_6_in( ArrayRowModule_3_io_V_wire_out_358 ),
       .io_VwirePorts_3_22_6_en( T1462 ),
       .io_VwirePorts_3_22_6_out( VwireModule_io_VwirePorts_3_22_6_out ),
       .io_VwirePorts_3_22_5_in( ArrayRowModule_3_io_V_wire_out_357 ),
       .io_VwirePorts_3_22_5_en( T1461 ),
       .io_VwirePorts_3_22_5_out( VwireModule_io_VwirePorts_3_22_5_out ),
       .io_VwirePorts_3_22_4_in( ArrayRowModule_3_io_V_wire_out_356 ),
       .io_VwirePorts_3_22_4_en( T1460 ),
       .io_VwirePorts_3_22_4_out( VwireModule_io_VwirePorts_3_22_4_out ),
       .io_VwirePorts_3_22_3_in( ArrayRowModule_3_io_V_wire_out_355 ),
       .io_VwirePorts_3_22_3_en( T1459 ),
       .io_VwirePorts_3_22_3_out( VwireModule_io_VwirePorts_3_22_3_out ),
       .io_VwirePorts_3_22_2_in( ArrayRowModule_3_io_V_wire_out_354 ),
       .io_VwirePorts_3_22_2_en( T1458 ),
       .io_VwirePorts_3_22_2_out( VwireModule_io_VwirePorts_3_22_2_out ),
       .io_VwirePorts_3_22_1_in( ArrayRowModule_3_io_V_wire_out_353 ),
       .io_VwirePorts_3_22_1_en( T1457 ),
       .io_VwirePorts_3_22_1_out( VwireModule_io_VwirePorts_3_22_1_out ),
       .io_VwirePorts_3_22_0_in( ArrayRowModule_3_io_V_wire_out_352 ),
       .io_VwirePorts_3_22_0_en( T1456 ),
       .io_VwirePorts_3_22_0_out( VwireModule_io_VwirePorts_3_22_0_out ),
       .io_VwirePorts_3_21_15_in( ArrayRowModule_3_io_V_wire_out_351 ),
       .io_VwirePorts_3_21_15_en( T1455 ),
       .io_VwirePorts_3_21_15_out( VwireModule_io_VwirePorts_3_21_15_out ),
       .io_VwirePorts_3_21_14_in( ArrayRowModule_3_io_V_wire_out_350 ),
       .io_VwirePorts_3_21_14_en( T1454 ),
       .io_VwirePorts_3_21_14_out( VwireModule_io_VwirePorts_3_21_14_out ),
       .io_VwirePorts_3_21_13_in( ArrayRowModule_3_io_V_wire_out_349 ),
       .io_VwirePorts_3_21_13_en( T1453 ),
       .io_VwirePorts_3_21_13_out( VwireModule_io_VwirePorts_3_21_13_out ),
       .io_VwirePorts_3_21_12_in( ArrayRowModule_3_io_V_wire_out_348 ),
       .io_VwirePorts_3_21_12_en( T1452 ),
       .io_VwirePorts_3_21_12_out( VwireModule_io_VwirePorts_3_21_12_out ),
       .io_VwirePorts_3_21_11_in( ArrayRowModule_3_io_V_wire_out_347 ),
       .io_VwirePorts_3_21_11_en( T1451 ),
       .io_VwirePorts_3_21_11_out( VwireModule_io_VwirePorts_3_21_11_out ),
       .io_VwirePorts_3_21_10_in( ArrayRowModule_3_io_V_wire_out_346 ),
       .io_VwirePorts_3_21_10_en( T1450 ),
       .io_VwirePorts_3_21_10_out( VwireModule_io_VwirePorts_3_21_10_out ),
       .io_VwirePorts_3_21_9_in( ArrayRowModule_3_io_V_wire_out_345 ),
       .io_VwirePorts_3_21_9_en( T1449 ),
       .io_VwirePorts_3_21_9_out( VwireModule_io_VwirePorts_3_21_9_out ),
       .io_VwirePorts_3_21_8_in( ArrayRowModule_3_io_V_wire_out_344 ),
       .io_VwirePorts_3_21_8_en( T1448 ),
       .io_VwirePorts_3_21_8_out( VwireModule_io_VwirePorts_3_21_8_out ),
       .io_VwirePorts_3_21_7_in( ArrayRowModule_3_io_V_wire_out_343 ),
       .io_VwirePorts_3_21_7_en( T1447 ),
       .io_VwirePorts_3_21_7_out( VwireModule_io_VwirePorts_3_21_7_out ),
       .io_VwirePorts_3_21_6_in( ArrayRowModule_3_io_V_wire_out_342 ),
       .io_VwirePorts_3_21_6_en( T1446 ),
       .io_VwirePorts_3_21_6_out( VwireModule_io_VwirePorts_3_21_6_out ),
       .io_VwirePorts_3_21_5_in( ArrayRowModule_3_io_V_wire_out_341 ),
       .io_VwirePorts_3_21_5_en( T1445 ),
       .io_VwirePorts_3_21_5_out( VwireModule_io_VwirePorts_3_21_5_out ),
       .io_VwirePorts_3_21_4_in( ArrayRowModule_3_io_V_wire_out_340 ),
       .io_VwirePorts_3_21_4_en( T1444 ),
       .io_VwirePorts_3_21_4_out( VwireModule_io_VwirePorts_3_21_4_out ),
       .io_VwirePorts_3_21_3_in( ArrayRowModule_3_io_V_wire_out_339 ),
       .io_VwirePorts_3_21_3_en( T1443 ),
       .io_VwirePorts_3_21_3_out( VwireModule_io_VwirePorts_3_21_3_out ),
       .io_VwirePorts_3_21_2_in( ArrayRowModule_3_io_V_wire_out_338 ),
       .io_VwirePorts_3_21_2_en( T1442 ),
       .io_VwirePorts_3_21_2_out( VwireModule_io_VwirePorts_3_21_2_out ),
       .io_VwirePorts_3_21_1_in( ArrayRowModule_3_io_V_wire_out_337 ),
       .io_VwirePorts_3_21_1_en( T1441 ),
       .io_VwirePorts_3_21_1_out( VwireModule_io_VwirePorts_3_21_1_out ),
       .io_VwirePorts_3_21_0_in( ArrayRowModule_3_io_V_wire_out_336 ),
       .io_VwirePorts_3_21_0_en( T1440 ),
       .io_VwirePorts_3_21_0_out( VwireModule_io_VwirePorts_3_21_0_out ),
       .io_VwirePorts_3_20_15_in( ArrayRowModule_3_io_V_wire_out_335 ),
       .io_VwirePorts_3_20_15_en( T1439 ),
       .io_VwirePorts_3_20_15_out( VwireModule_io_VwirePorts_3_20_15_out ),
       .io_VwirePorts_3_20_14_in( ArrayRowModule_3_io_V_wire_out_334 ),
       .io_VwirePorts_3_20_14_en( T1438 ),
       .io_VwirePorts_3_20_14_out( VwireModule_io_VwirePorts_3_20_14_out ),
       .io_VwirePorts_3_20_13_in( ArrayRowModule_3_io_V_wire_out_333 ),
       .io_VwirePorts_3_20_13_en( T1437 ),
       .io_VwirePorts_3_20_13_out( VwireModule_io_VwirePorts_3_20_13_out ),
       .io_VwirePorts_3_20_12_in( ArrayRowModule_3_io_V_wire_out_332 ),
       .io_VwirePorts_3_20_12_en( T1436 ),
       .io_VwirePorts_3_20_12_out( VwireModule_io_VwirePorts_3_20_12_out ),
       .io_VwirePorts_3_20_11_in( ArrayRowModule_3_io_V_wire_out_331 ),
       .io_VwirePorts_3_20_11_en( T1435 ),
       .io_VwirePorts_3_20_11_out( VwireModule_io_VwirePorts_3_20_11_out ),
       .io_VwirePorts_3_20_10_in( ArrayRowModule_3_io_V_wire_out_330 ),
       .io_VwirePorts_3_20_10_en( T1434 ),
       .io_VwirePorts_3_20_10_out( VwireModule_io_VwirePorts_3_20_10_out ),
       .io_VwirePorts_3_20_9_in( ArrayRowModule_3_io_V_wire_out_329 ),
       .io_VwirePorts_3_20_9_en( T1433 ),
       .io_VwirePorts_3_20_9_out( VwireModule_io_VwirePorts_3_20_9_out ),
       .io_VwirePorts_3_20_8_in( ArrayRowModule_3_io_V_wire_out_328 ),
       .io_VwirePorts_3_20_8_en( T1432 ),
       .io_VwirePorts_3_20_8_out( VwireModule_io_VwirePorts_3_20_8_out ),
       .io_VwirePorts_3_20_7_in( ArrayRowModule_3_io_V_wire_out_327 ),
       .io_VwirePorts_3_20_7_en( T1431 ),
       .io_VwirePorts_3_20_7_out( VwireModule_io_VwirePorts_3_20_7_out ),
       .io_VwirePorts_3_20_6_in( ArrayRowModule_3_io_V_wire_out_326 ),
       .io_VwirePorts_3_20_6_en( T1430 ),
       .io_VwirePorts_3_20_6_out( VwireModule_io_VwirePorts_3_20_6_out ),
       .io_VwirePorts_3_20_5_in( ArrayRowModule_3_io_V_wire_out_325 ),
       .io_VwirePorts_3_20_5_en( T1429 ),
       .io_VwirePorts_3_20_5_out( VwireModule_io_VwirePorts_3_20_5_out ),
       .io_VwirePorts_3_20_4_in( ArrayRowModule_3_io_V_wire_out_324 ),
       .io_VwirePorts_3_20_4_en( T1428 ),
       .io_VwirePorts_3_20_4_out( VwireModule_io_VwirePorts_3_20_4_out ),
       .io_VwirePorts_3_20_3_in( ArrayRowModule_3_io_V_wire_out_323 ),
       .io_VwirePorts_3_20_3_en( T1427 ),
       .io_VwirePorts_3_20_3_out( VwireModule_io_VwirePorts_3_20_3_out ),
       .io_VwirePorts_3_20_2_in( ArrayRowModule_3_io_V_wire_out_322 ),
       .io_VwirePorts_3_20_2_en( T1426 ),
       .io_VwirePorts_3_20_2_out( VwireModule_io_VwirePorts_3_20_2_out ),
       .io_VwirePorts_3_20_1_in( ArrayRowModule_3_io_V_wire_out_321 ),
       .io_VwirePorts_3_20_1_en( T1425 ),
       .io_VwirePorts_3_20_1_out( VwireModule_io_VwirePorts_3_20_1_out ),
       .io_VwirePorts_3_20_0_in( ArrayRowModule_3_io_V_wire_out_320 ),
       .io_VwirePorts_3_20_0_en( T1424 ),
       .io_VwirePorts_3_20_0_out( VwireModule_io_VwirePorts_3_20_0_out ),
       .io_VwirePorts_3_19_15_in( ArrayRowModule_3_io_V_wire_out_319 ),
       .io_VwirePorts_3_19_15_en( T1423 ),
       .io_VwirePorts_3_19_15_out( VwireModule_io_VwirePorts_3_19_15_out ),
       .io_VwirePorts_3_19_14_in( ArrayRowModule_3_io_V_wire_out_318 ),
       .io_VwirePorts_3_19_14_en( T1422 ),
       .io_VwirePorts_3_19_14_out( VwireModule_io_VwirePorts_3_19_14_out ),
       .io_VwirePorts_3_19_13_in( ArrayRowModule_3_io_V_wire_out_317 ),
       .io_VwirePorts_3_19_13_en( T1421 ),
       .io_VwirePorts_3_19_13_out( VwireModule_io_VwirePorts_3_19_13_out ),
       .io_VwirePorts_3_19_12_in( ArrayRowModule_3_io_V_wire_out_316 ),
       .io_VwirePorts_3_19_12_en( T1420 ),
       .io_VwirePorts_3_19_12_out( VwireModule_io_VwirePorts_3_19_12_out ),
       .io_VwirePorts_3_19_11_in( ArrayRowModule_3_io_V_wire_out_315 ),
       .io_VwirePorts_3_19_11_en( T1419 ),
       .io_VwirePorts_3_19_11_out( VwireModule_io_VwirePorts_3_19_11_out ),
       .io_VwirePorts_3_19_10_in( ArrayRowModule_3_io_V_wire_out_314 ),
       .io_VwirePorts_3_19_10_en( T1418 ),
       .io_VwirePorts_3_19_10_out( VwireModule_io_VwirePorts_3_19_10_out ),
       .io_VwirePorts_3_19_9_in( ArrayRowModule_3_io_V_wire_out_313 ),
       .io_VwirePorts_3_19_9_en( T1417 ),
       .io_VwirePorts_3_19_9_out( VwireModule_io_VwirePorts_3_19_9_out ),
       .io_VwirePorts_3_19_8_in( ArrayRowModule_3_io_V_wire_out_312 ),
       .io_VwirePorts_3_19_8_en( T1416 ),
       .io_VwirePorts_3_19_8_out( VwireModule_io_VwirePorts_3_19_8_out ),
       .io_VwirePorts_3_19_7_in( ArrayRowModule_3_io_V_wire_out_311 ),
       .io_VwirePorts_3_19_7_en( T1415 ),
       .io_VwirePorts_3_19_7_out( VwireModule_io_VwirePorts_3_19_7_out ),
       .io_VwirePorts_3_19_6_in( ArrayRowModule_3_io_V_wire_out_310 ),
       .io_VwirePorts_3_19_6_en( T1414 ),
       .io_VwirePorts_3_19_6_out( VwireModule_io_VwirePorts_3_19_6_out ),
       .io_VwirePorts_3_19_5_in( ArrayRowModule_3_io_V_wire_out_309 ),
       .io_VwirePorts_3_19_5_en( T1413 ),
       .io_VwirePorts_3_19_5_out( VwireModule_io_VwirePorts_3_19_5_out ),
       .io_VwirePorts_3_19_4_in( ArrayRowModule_3_io_V_wire_out_308 ),
       .io_VwirePorts_3_19_4_en( T1412 ),
       .io_VwirePorts_3_19_4_out( VwireModule_io_VwirePorts_3_19_4_out ),
       .io_VwirePorts_3_19_3_in( ArrayRowModule_3_io_V_wire_out_307 ),
       .io_VwirePorts_3_19_3_en( T1411 ),
       .io_VwirePorts_3_19_3_out( VwireModule_io_VwirePorts_3_19_3_out ),
       .io_VwirePorts_3_19_2_in( ArrayRowModule_3_io_V_wire_out_306 ),
       .io_VwirePorts_3_19_2_en( T1410 ),
       .io_VwirePorts_3_19_2_out( VwireModule_io_VwirePorts_3_19_2_out ),
       .io_VwirePorts_3_19_1_in( ArrayRowModule_3_io_V_wire_out_305 ),
       .io_VwirePorts_3_19_1_en( T1409 ),
       .io_VwirePorts_3_19_1_out( VwireModule_io_VwirePorts_3_19_1_out ),
       .io_VwirePorts_3_19_0_in( ArrayRowModule_3_io_V_wire_out_304 ),
       .io_VwirePorts_3_19_0_en( T1408 ),
       .io_VwirePorts_3_19_0_out( VwireModule_io_VwirePorts_3_19_0_out ),
       .io_VwirePorts_3_18_15_in( ArrayRowModule_3_io_V_wire_out_303 ),
       .io_VwirePorts_3_18_15_en( T1407 ),
       .io_VwirePorts_3_18_15_out( VwireModule_io_VwirePorts_3_18_15_out ),
       .io_VwirePorts_3_18_14_in( ArrayRowModule_3_io_V_wire_out_302 ),
       .io_VwirePorts_3_18_14_en( T1406 ),
       .io_VwirePorts_3_18_14_out( VwireModule_io_VwirePorts_3_18_14_out ),
       .io_VwirePorts_3_18_13_in( ArrayRowModule_3_io_V_wire_out_301 ),
       .io_VwirePorts_3_18_13_en( T1405 ),
       .io_VwirePorts_3_18_13_out( VwireModule_io_VwirePorts_3_18_13_out ),
       .io_VwirePorts_3_18_12_in( ArrayRowModule_3_io_V_wire_out_300 ),
       .io_VwirePorts_3_18_12_en( T1404 ),
       .io_VwirePorts_3_18_12_out( VwireModule_io_VwirePorts_3_18_12_out ),
       .io_VwirePorts_3_18_11_in( ArrayRowModule_3_io_V_wire_out_299 ),
       .io_VwirePorts_3_18_11_en( T1403 ),
       .io_VwirePorts_3_18_11_out( VwireModule_io_VwirePorts_3_18_11_out ),
       .io_VwirePorts_3_18_10_in( ArrayRowModule_3_io_V_wire_out_298 ),
       .io_VwirePorts_3_18_10_en( T1402 ),
       .io_VwirePorts_3_18_10_out( VwireModule_io_VwirePorts_3_18_10_out ),
       .io_VwirePorts_3_18_9_in( ArrayRowModule_3_io_V_wire_out_297 ),
       .io_VwirePorts_3_18_9_en( T1401 ),
       .io_VwirePorts_3_18_9_out( VwireModule_io_VwirePorts_3_18_9_out ),
       .io_VwirePorts_3_18_8_in( ArrayRowModule_3_io_V_wire_out_296 ),
       .io_VwirePorts_3_18_8_en( T1400 ),
       .io_VwirePorts_3_18_8_out( VwireModule_io_VwirePorts_3_18_8_out ),
       .io_VwirePorts_3_18_7_in( ArrayRowModule_3_io_V_wire_out_295 ),
       .io_VwirePorts_3_18_7_en( T1399 ),
       .io_VwirePorts_3_18_7_out( VwireModule_io_VwirePorts_3_18_7_out ),
       .io_VwirePorts_3_18_6_in( ArrayRowModule_3_io_V_wire_out_294 ),
       .io_VwirePorts_3_18_6_en( T1398 ),
       .io_VwirePorts_3_18_6_out( VwireModule_io_VwirePorts_3_18_6_out ),
       .io_VwirePorts_3_18_5_in( ArrayRowModule_3_io_V_wire_out_293 ),
       .io_VwirePorts_3_18_5_en( T1397 ),
       .io_VwirePorts_3_18_5_out( VwireModule_io_VwirePorts_3_18_5_out ),
       .io_VwirePorts_3_18_4_in( ArrayRowModule_3_io_V_wire_out_292 ),
       .io_VwirePorts_3_18_4_en( T1396 ),
       .io_VwirePorts_3_18_4_out( VwireModule_io_VwirePorts_3_18_4_out ),
       .io_VwirePorts_3_18_3_in( ArrayRowModule_3_io_V_wire_out_291 ),
       .io_VwirePorts_3_18_3_en( T1395 ),
       .io_VwirePorts_3_18_3_out( VwireModule_io_VwirePorts_3_18_3_out ),
       .io_VwirePorts_3_18_2_in( ArrayRowModule_3_io_V_wire_out_290 ),
       .io_VwirePorts_3_18_2_en( T1394 ),
       .io_VwirePorts_3_18_2_out( VwireModule_io_VwirePorts_3_18_2_out ),
       .io_VwirePorts_3_18_1_in( ArrayRowModule_3_io_V_wire_out_289 ),
       .io_VwirePorts_3_18_1_en( T1393 ),
       .io_VwirePorts_3_18_1_out( VwireModule_io_VwirePorts_3_18_1_out ),
       .io_VwirePorts_3_18_0_in( ArrayRowModule_3_io_V_wire_out_288 ),
       .io_VwirePorts_3_18_0_en( T1392 ),
       .io_VwirePorts_3_18_0_out( VwireModule_io_VwirePorts_3_18_0_out ),
       .io_VwirePorts_3_17_15_in( ArrayRowModule_3_io_V_wire_out_287 ),
       .io_VwirePorts_3_17_15_en( T1391 ),
       .io_VwirePorts_3_17_15_out( VwireModule_io_VwirePorts_3_17_15_out ),
       .io_VwirePorts_3_17_14_in( ArrayRowModule_3_io_V_wire_out_286 ),
       .io_VwirePorts_3_17_14_en( T1390 ),
       .io_VwirePorts_3_17_14_out( VwireModule_io_VwirePorts_3_17_14_out ),
       .io_VwirePorts_3_17_13_in( ArrayRowModule_3_io_V_wire_out_285 ),
       .io_VwirePorts_3_17_13_en( T1389 ),
       .io_VwirePorts_3_17_13_out( VwireModule_io_VwirePorts_3_17_13_out ),
       .io_VwirePorts_3_17_12_in( ArrayRowModule_3_io_V_wire_out_284 ),
       .io_VwirePorts_3_17_12_en( T1388 ),
       .io_VwirePorts_3_17_12_out( VwireModule_io_VwirePorts_3_17_12_out ),
       .io_VwirePorts_3_17_11_in( ArrayRowModule_3_io_V_wire_out_283 ),
       .io_VwirePorts_3_17_11_en( T1387 ),
       .io_VwirePorts_3_17_11_out( VwireModule_io_VwirePorts_3_17_11_out ),
       .io_VwirePorts_3_17_10_in( ArrayRowModule_3_io_V_wire_out_282 ),
       .io_VwirePorts_3_17_10_en( T1386 ),
       .io_VwirePorts_3_17_10_out( VwireModule_io_VwirePorts_3_17_10_out ),
       .io_VwirePorts_3_17_9_in( ArrayRowModule_3_io_V_wire_out_281 ),
       .io_VwirePorts_3_17_9_en( T1385 ),
       .io_VwirePorts_3_17_9_out( VwireModule_io_VwirePorts_3_17_9_out ),
       .io_VwirePorts_3_17_8_in( ArrayRowModule_3_io_V_wire_out_280 ),
       .io_VwirePorts_3_17_8_en( T1384 ),
       .io_VwirePorts_3_17_8_out( VwireModule_io_VwirePorts_3_17_8_out ),
       .io_VwirePorts_3_17_7_in( ArrayRowModule_3_io_V_wire_out_279 ),
       .io_VwirePorts_3_17_7_en( T1383 ),
       .io_VwirePorts_3_17_7_out( VwireModule_io_VwirePorts_3_17_7_out ),
       .io_VwirePorts_3_17_6_in( ArrayRowModule_3_io_V_wire_out_278 ),
       .io_VwirePorts_3_17_6_en( T1382 ),
       .io_VwirePorts_3_17_6_out( VwireModule_io_VwirePorts_3_17_6_out ),
       .io_VwirePorts_3_17_5_in( ArrayRowModule_3_io_V_wire_out_277 ),
       .io_VwirePorts_3_17_5_en( T1381 ),
       .io_VwirePorts_3_17_5_out( VwireModule_io_VwirePorts_3_17_5_out ),
       .io_VwirePorts_3_17_4_in( ArrayRowModule_3_io_V_wire_out_276 ),
       .io_VwirePorts_3_17_4_en( T1380 ),
       .io_VwirePorts_3_17_4_out( VwireModule_io_VwirePorts_3_17_4_out ),
       .io_VwirePorts_3_17_3_in( ArrayRowModule_3_io_V_wire_out_275 ),
       .io_VwirePorts_3_17_3_en( T1379 ),
       .io_VwirePorts_3_17_3_out( VwireModule_io_VwirePorts_3_17_3_out ),
       .io_VwirePorts_3_17_2_in( ArrayRowModule_3_io_V_wire_out_274 ),
       .io_VwirePorts_3_17_2_en( T1378 ),
       .io_VwirePorts_3_17_2_out( VwireModule_io_VwirePorts_3_17_2_out ),
       .io_VwirePorts_3_17_1_in( ArrayRowModule_3_io_V_wire_out_273 ),
       .io_VwirePorts_3_17_1_en( T1377 ),
       .io_VwirePorts_3_17_1_out( VwireModule_io_VwirePorts_3_17_1_out ),
       .io_VwirePorts_3_17_0_in( ArrayRowModule_3_io_V_wire_out_272 ),
       .io_VwirePorts_3_17_0_en( T1376 ),
       .io_VwirePorts_3_17_0_out( VwireModule_io_VwirePorts_3_17_0_out ),
       .io_VwirePorts_3_16_15_in( ArrayRowModule_3_io_V_wire_out_271 ),
       .io_VwirePorts_3_16_15_en( T1375 ),
       .io_VwirePorts_3_16_15_out( VwireModule_io_VwirePorts_3_16_15_out ),
       .io_VwirePorts_3_16_14_in( ArrayRowModule_3_io_V_wire_out_270 ),
       .io_VwirePorts_3_16_14_en( T1374 ),
       .io_VwirePorts_3_16_14_out( VwireModule_io_VwirePorts_3_16_14_out ),
       .io_VwirePorts_3_16_13_in( ArrayRowModule_3_io_V_wire_out_269 ),
       .io_VwirePorts_3_16_13_en( T1373 ),
       .io_VwirePorts_3_16_13_out( VwireModule_io_VwirePorts_3_16_13_out ),
       .io_VwirePorts_3_16_12_in( ArrayRowModule_3_io_V_wire_out_268 ),
       .io_VwirePorts_3_16_12_en( T1372 ),
       .io_VwirePorts_3_16_12_out( VwireModule_io_VwirePorts_3_16_12_out ),
       .io_VwirePorts_3_16_11_in( ArrayRowModule_3_io_V_wire_out_267 ),
       .io_VwirePorts_3_16_11_en( T1371 ),
       .io_VwirePorts_3_16_11_out( VwireModule_io_VwirePorts_3_16_11_out ),
       .io_VwirePorts_3_16_10_in( ArrayRowModule_3_io_V_wire_out_266 ),
       .io_VwirePorts_3_16_10_en( T1370 ),
       .io_VwirePorts_3_16_10_out( VwireModule_io_VwirePorts_3_16_10_out ),
       .io_VwirePorts_3_16_9_in( ArrayRowModule_3_io_V_wire_out_265 ),
       .io_VwirePorts_3_16_9_en( T1369 ),
       .io_VwirePorts_3_16_9_out( VwireModule_io_VwirePorts_3_16_9_out ),
       .io_VwirePorts_3_16_8_in( ArrayRowModule_3_io_V_wire_out_264 ),
       .io_VwirePorts_3_16_8_en( T1368 ),
       .io_VwirePorts_3_16_8_out( VwireModule_io_VwirePorts_3_16_8_out ),
       .io_VwirePorts_3_16_7_in( ArrayRowModule_3_io_V_wire_out_263 ),
       .io_VwirePorts_3_16_7_en( T1367 ),
       .io_VwirePorts_3_16_7_out( VwireModule_io_VwirePorts_3_16_7_out ),
       .io_VwirePorts_3_16_6_in( ArrayRowModule_3_io_V_wire_out_262 ),
       .io_VwirePorts_3_16_6_en( T1366 ),
       .io_VwirePorts_3_16_6_out( VwireModule_io_VwirePorts_3_16_6_out ),
       .io_VwirePorts_3_16_5_in( ArrayRowModule_3_io_V_wire_out_261 ),
       .io_VwirePorts_3_16_5_en( T1365 ),
       .io_VwirePorts_3_16_5_out( VwireModule_io_VwirePorts_3_16_5_out ),
       .io_VwirePorts_3_16_4_in( ArrayRowModule_3_io_V_wire_out_260 ),
       .io_VwirePorts_3_16_4_en( T1364 ),
       .io_VwirePorts_3_16_4_out( VwireModule_io_VwirePorts_3_16_4_out ),
       .io_VwirePorts_3_16_3_in( ArrayRowModule_3_io_V_wire_out_259 ),
       .io_VwirePorts_3_16_3_en( T1363 ),
       .io_VwirePorts_3_16_3_out( VwireModule_io_VwirePorts_3_16_3_out ),
       .io_VwirePorts_3_16_2_in( ArrayRowModule_3_io_V_wire_out_258 ),
       .io_VwirePorts_3_16_2_en( T1362 ),
       .io_VwirePorts_3_16_2_out( VwireModule_io_VwirePorts_3_16_2_out ),
       .io_VwirePorts_3_16_1_in( ArrayRowModule_3_io_V_wire_out_257 ),
       .io_VwirePorts_3_16_1_en( T1361 ),
       .io_VwirePorts_3_16_1_out( VwireModule_io_VwirePorts_3_16_1_out ),
       .io_VwirePorts_3_16_0_in( ArrayRowModule_3_io_V_wire_out_256 ),
       .io_VwirePorts_3_16_0_en( T1360 ),
       .io_VwirePorts_3_16_0_out( VwireModule_io_VwirePorts_3_16_0_out ),
       .io_VwirePorts_3_15_15_in( ArrayRowModule_3_io_V_wire_out_255 ),
       .io_VwirePorts_3_15_15_en( T1359 ),
       .io_VwirePorts_3_15_15_out( VwireModule_io_VwirePorts_3_15_15_out ),
       .io_VwirePorts_3_15_14_in( ArrayRowModule_3_io_V_wire_out_254 ),
       .io_VwirePorts_3_15_14_en( T1358 ),
       .io_VwirePorts_3_15_14_out( VwireModule_io_VwirePorts_3_15_14_out ),
       .io_VwirePorts_3_15_13_in( ArrayRowModule_3_io_V_wire_out_253 ),
       .io_VwirePorts_3_15_13_en( T1357 ),
       .io_VwirePorts_3_15_13_out( VwireModule_io_VwirePorts_3_15_13_out ),
       .io_VwirePorts_3_15_12_in( ArrayRowModule_3_io_V_wire_out_252 ),
       .io_VwirePorts_3_15_12_en( T1356 ),
       .io_VwirePorts_3_15_12_out( VwireModule_io_VwirePorts_3_15_12_out ),
       .io_VwirePorts_3_15_11_in( ArrayRowModule_3_io_V_wire_out_251 ),
       .io_VwirePorts_3_15_11_en( T1355 ),
       .io_VwirePorts_3_15_11_out( VwireModule_io_VwirePorts_3_15_11_out ),
       .io_VwirePorts_3_15_10_in( ArrayRowModule_3_io_V_wire_out_250 ),
       .io_VwirePorts_3_15_10_en( T1354 ),
       .io_VwirePorts_3_15_10_out( VwireModule_io_VwirePorts_3_15_10_out ),
       .io_VwirePorts_3_15_9_in( ArrayRowModule_3_io_V_wire_out_249 ),
       .io_VwirePorts_3_15_9_en( T1353 ),
       .io_VwirePorts_3_15_9_out( VwireModule_io_VwirePorts_3_15_9_out ),
       .io_VwirePorts_3_15_8_in( ArrayRowModule_3_io_V_wire_out_248 ),
       .io_VwirePorts_3_15_8_en( T1352 ),
       .io_VwirePorts_3_15_8_out( VwireModule_io_VwirePorts_3_15_8_out ),
       .io_VwirePorts_3_15_7_in( ArrayRowModule_3_io_V_wire_out_247 ),
       .io_VwirePorts_3_15_7_en( T1351 ),
       .io_VwirePorts_3_15_7_out( VwireModule_io_VwirePorts_3_15_7_out ),
       .io_VwirePorts_3_15_6_in( ArrayRowModule_3_io_V_wire_out_246 ),
       .io_VwirePorts_3_15_6_en( T1350 ),
       .io_VwirePorts_3_15_6_out( VwireModule_io_VwirePorts_3_15_6_out ),
       .io_VwirePorts_3_15_5_in( ArrayRowModule_3_io_V_wire_out_245 ),
       .io_VwirePorts_3_15_5_en( T1349 ),
       .io_VwirePorts_3_15_5_out( VwireModule_io_VwirePorts_3_15_5_out ),
       .io_VwirePorts_3_15_4_in( ArrayRowModule_3_io_V_wire_out_244 ),
       .io_VwirePorts_3_15_4_en( T1348 ),
       .io_VwirePorts_3_15_4_out( VwireModule_io_VwirePorts_3_15_4_out ),
       .io_VwirePorts_3_15_3_in( ArrayRowModule_3_io_V_wire_out_243 ),
       .io_VwirePorts_3_15_3_en( T1347 ),
       .io_VwirePorts_3_15_3_out( VwireModule_io_VwirePorts_3_15_3_out ),
       .io_VwirePorts_3_15_2_in( ArrayRowModule_3_io_V_wire_out_242 ),
       .io_VwirePorts_3_15_2_en( T1346 ),
       .io_VwirePorts_3_15_2_out( VwireModule_io_VwirePorts_3_15_2_out ),
       .io_VwirePorts_3_15_1_in( ArrayRowModule_3_io_V_wire_out_241 ),
       .io_VwirePorts_3_15_1_en( T1345 ),
       .io_VwirePorts_3_15_1_out( VwireModule_io_VwirePorts_3_15_1_out ),
       .io_VwirePorts_3_15_0_in( ArrayRowModule_3_io_V_wire_out_240 ),
       .io_VwirePorts_3_15_0_en( T1344 ),
       .io_VwirePorts_3_15_0_out( VwireModule_io_VwirePorts_3_15_0_out ),
       .io_VwirePorts_3_14_15_in( ArrayRowModule_3_io_V_wire_out_239 ),
       .io_VwirePorts_3_14_15_en( T1343 ),
       .io_VwirePorts_3_14_15_out( VwireModule_io_VwirePorts_3_14_15_out ),
       .io_VwirePorts_3_14_14_in( ArrayRowModule_3_io_V_wire_out_238 ),
       .io_VwirePorts_3_14_14_en( T1342 ),
       .io_VwirePorts_3_14_14_out( VwireModule_io_VwirePorts_3_14_14_out ),
       .io_VwirePorts_3_14_13_in( ArrayRowModule_3_io_V_wire_out_237 ),
       .io_VwirePorts_3_14_13_en( T1341 ),
       .io_VwirePorts_3_14_13_out( VwireModule_io_VwirePorts_3_14_13_out ),
       .io_VwirePorts_3_14_12_in( ArrayRowModule_3_io_V_wire_out_236 ),
       .io_VwirePorts_3_14_12_en( T1340 ),
       .io_VwirePorts_3_14_12_out( VwireModule_io_VwirePorts_3_14_12_out ),
       .io_VwirePorts_3_14_11_in( ArrayRowModule_3_io_V_wire_out_235 ),
       .io_VwirePorts_3_14_11_en( T1339 ),
       .io_VwirePorts_3_14_11_out( VwireModule_io_VwirePorts_3_14_11_out ),
       .io_VwirePorts_3_14_10_in( ArrayRowModule_3_io_V_wire_out_234 ),
       .io_VwirePorts_3_14_10_en( T1338 ),
       .io_VwirePorts_3_14_10_out( VwireModule_io_VwirePorts_3_14_10_out ),
       .io_VwirePorts_3_14_9_in( ArrayRowModule_3_io_V_wire_out_233 ),
       .io_VwirePorts_3_14_9_en( T1337 ),
       .io_VwirePorts_3_14_9_out( VwireModule_io_VwirePorts_3_14_9_out ),
       .io_VwirePorts_3_14_8_in( ArrayRowModule_3_io_V_wire_out_232 ),
       .io_VwirePorts_3_14_8_en( T1336 ),
       .io_VwirePorts_3_14_8_out( VwireModule_io_VwirePorts_3_14_8_out ),
       .io_VwirePorts_3_14_7_in( ArrayRowModule_3_io_V_wire_out_231 ),
       .io_VwirePorts_3_14_7_en( T1335 ),
       .io_VwirePorts_3_14_7_out( VwireModule_io_VwirePorts_3_14_7_out ),
       .io_VwirePorts_3_14_6_in( ArrayRowModule_3_io_V_wire_out_230 ),
       .io_VwirePorts_3_14_6_en( T1334 ),
       .io_VwirePorts_3_14_6_out( VwireModule_io_VwirePorts_3_14_6_out ),
       .io_VwirePorts_3_14_5_in( ArrayRowModule_3_io_V_wire_out_229 ),
       .io_VwirePorts_3_14_5_en( T1333 ),
       .io_VwirePorts_3_14_5_out( VwireModule_io_VwirePorts_3_14_5_out ),
       .io_VwirePorts_3_14_4_in( ArrayRowModule_3_io_V_wire_out_228 ),
       .io_VwirePorts_3_14_4_en( T1332 ),
       .io_VwirePorts_3_14_4_out( VwireModule_io_VwirePorts_3_14_4_out ),
       .io_VwirePorts_3_14_3_in( ArrayRowModule_3_io_V_wire_out_227 ),
       .io_VwirePorts_3_14_3_en( T1331 ),
       .io_VwirePorts_3_14_3_out( VwireModule_io_VwirePorts_3_14_3_out ),
       .io_VwirePorts_3_14_2_in( ArrayRowModule_3_io_V_wire_out_226 ),
       .io_VwirePorts_3_14_2_en( T1330 ),
       .io_VwirePorts_3_14_2_out( VwireModule_io_VwirePorts_3_14_2_out ),
       .io_VwirePorts_3_14_1_in( ArrayRowModule_3_io_V_wire_out_225 ),
       .io_VwirePorts_3_14_1_en( T1329 ),
       .io_VwirePorts_3_14_1_out( VwireModule_io_VwirePorts_3_14_1_out ),
       .io_VwirePorts_3_14_0_in( ArrayRowModule_3_io_V_wire_out_224 ),
       .io_VwirePorts_3_14_0_en( T1328 ),
       .io_VwirePorts_3_14_0_out( VwireModule_io_VwirePorts_3_14_0_out ),
       .io_VwirePorts_3_13_15_in( ArrayRowModule_3_io_V_wire_out_223 ),
       .io_VwirePorts_3_13_15_en( T1327 ),
       .io_VwirePorts_3_13_15_out( VwireModule_io_VwirePorts_3_13_15_out ),
       .io_VwirePorts_3_13_14_in( ArrayRowModule_3_io_V_wire_out_222 ),
       .io_VwirePorts_3_13_14_en( T1326 ),
       .io_VwirePorts_3_13_14_out( VwireModule_io_VwirePorts_3_13_14_out ),
       .io_VwirePorts_3_13_13_in( ArrayRowModule_3_io_V_wire_out_221 ),
       .io_VwirePorts_3_13_13_en( T1325 ),
       .io_VwirePorts_3_13_13_out( VwireModule_io_VwirePorts_3_13_13_out ),
       .io_VwirePorts_3_13_12_in( ArrayRowModule_3_io_V_wire_out_220 ),
       .io_VwirePorts_3_13_12_en( T1324 ),
       .io_VwirePorts_3_13_12_out( VwireModule_io_VwirePorts_3_13_12_out ),
       .io_VwirePorts_3_13_11_in( ArrayRowModule_3_io_V_wire_out_219 ),
       .io_VwirePorts_3_13_11_en( T1323 ),
       .io_VwirePorts_3_13_11_out( VwireModule_io_VwirePorts_3_13_11_out ),
       .io_VwirePorts_3_13_10_in( ArrayRowModule_3_io_V_wire_out_218 ),
       .io_VwirePorts_3_13_10_en( T1322 ),
       .io_VwirePorts_3_13_10_out( VwireModule_io_VwirePorts_3_13_10_out ),
       .io_VwirePorts_3_13_9_in( ArrayRowModule_3_io_V_wire_out_217 ),
       .io_VwirePorts_3_13_9_en( T1321 ),
       .io_VwirePorts_3_13_9_out( VwireModule_io_VwirePorts_3_13_9_out ),
       .io_VwirePorts_3_13_8_in( ArrayRowModule_3_io_V_wire_out_216 ),
       .io_VwirePorts_3_13_8_en( T1320 ),
       .io_VwirePorts_3_13_8_out( VwireModule_io_VwirePorts_3_13_8_out ),
       .io_VwirePorts_3_13_7_in( ArrayRowModule_3_io_V_wire_out_215 ),
       .io_VwirePorts_3_13_7_en( T1319 ),
       .io_VwirePorts_3_13_7_out( VwireModule_io_VwirePorts_3_13_7_out ),
       .io_VwirePorts_3_13_6_in( ArrayRowModule_3_io_V_wire_out_214 ),
       .io_VwirePorts_3_13_6_en( T1318 ),
       .io_VwirePorts_3_13_6_out( VwireModule_io_VwirePorts_3_13_6_out ),
       .io_VwirePorts_3_13_5_in( ArrayRowModule_3_io_V_wire_out_213 ),
       .io_VwirePorts_3_13_5_en( T1317 ),
       .io_VwirePorts_3_13_5_out( VwireModule_io_VwirePorts_3_13_5_out ),
       .io_VwirePorts_3_13_4_in( ArrayRowModule_3_io_V_wire_out_212 ),
       .io_VwirePorts_3_13_4_en( T1316 ),
       .io_VwirePorts_3_13_4_out( VwireModule_io_VwirePorts_3_13_4_out ),
       .io_VwirePorts_3_13_3_in( ArrayRowModule_3_io_V_wire_out_211 ),
       .io_VwirePorts_3_13_3_en( T1315 ),
       .io_VwirePorts_3_13_3_out( VwireModule_io_VwirePorts_3_13_3_out ),
       .io_VwirePorts_3_13_2_in( ArrayRowModule_3_io_V_wire_out_210 ),
       .io_VwirePorts_3_13_2_en( T1314 ),
       .io_VwirePorts_3_13_2_out( VwireModule_io_VwirePorts_3_13_2_out ),
       .io_VwirePorts_3_13_1_in( ArrayRowModule_3_io_V_wire_out_209 ),
       .io_VwirePorts_3_13_1_en( T1313 ),
       .io_VwirePorts_3_13_1_out( VwireModule_io_VwirePorts_3_13_1_out ),
       .io_VwirePorts_3_13_0_in( ArrayRowModule_3_io_V_wire_out_208 ),
       .io_VwirePorts_3_13_0_en( T1312 ),
       .io_VwirePorts_3_13_0_out( VwireModule_io_VwirePorts_3_13_0_out ),
       .io_VwirePorts_3_12_15_in( ArrayRowModule_3_io_V_wire_out_207 ),
       .io_VwirePorts_3_12_15_en( T1311 ),
       .io_VwirePorts_3_12_15_out( VwireModule_io_VwirePorts_3_12_15_out ),
       .io_VwirePorts_3_12_14_in( ArrayRowModule_3_io_V_wire_out_206 ),
       .io_VwirePorts_3_12_14_en( T1310 ),
       .io_VwirePorts_3_12_14_out( VwireModule_io_VwirePorts_3_12_14_out ),
       .io_VwirePorts_3_12_13_in( ArrayRowModule_3_io_V_wire_out_205 ),
       .io_VwirePorts_3_12_13_en( T1309 ),
       .io_VwirePorts_3_12_13_out( VwireModule_io_VwirePorts_3_12_13_out ),
       .io_VwirePorts_3_12_12_in( ArrayRowModule_3_io_V_wire_out_204 ),
       .io_VwirePorts_3_12_12_en( T1308 ),
       .io_VwirePorts_3_12_12_out( VwireModule_io_VwirePorts_3_12_12_out ),
       .io_VwirePorts_3_12_11_in( ArrayRowModule_3_io_V_wire_out_203 ),
       .io_VwirePorts_3_12_11_en( T1307 ),
       .io_VwirePorts_3_12_11_out( VwireModule_io_VwirePorts_3_12_11_out ),
       .io_VwirePorts_3_12_10_in( ArrayRowModule_3_io_V_wire_out_202 ),
       .io_VwirePorts_3_12_10_en( T1306 ),
       .io_VwirePorts_3_12_10_out( VwireModule_io_VwirePorts_3_12_10_out ),
       .io_VwirePorts_3_12_9_in( ArrayRowModule_3_io_V_wire_out_201 ),
       .io_VwirePorts_3_12_9_en( T1305 ),
       .io_VwirePorts_3_12_9_out( VwireModule_io_VwirePorts_3_12_9_out ),
       .io_VwirePorts_3_12_8_in( ArrayRowModule_3_io_V_wire_out_200 ),
       .io_VwirePorts_3_12_8_en( T1304 ),
       .io_VwirePorts_3_12_8_out( VwireModule_io_VwirePorts_3_12_8_out ),
       .io_VwirePorts_3_12_7_in( ArrayRowModule_3_io_V_wire_out_199 ),
       .io_VwirePorts_3_12_7_en( T1303 ),
       .io_VwirePorts_3_12_7_out( VwireModule_io_VwirePorts_3_12_7_out ),
       .io_VwirePorts_3_12_6_in( ArrayRowModule_3_io_V_wire_out_198 ),
       .io_VwirePorts_3_12_6_en( T1302 ),
       .io_VwirePorts_3_12_6_out( VwireModule_io_VwirePorts_3_12_6_out ),
       .io_VwirePorts_3_12_5_in( ArrayRowModule_3_io_V_wire_out_197 ),
       .io_VwirePorts_3_12_5_en( T1301 ),
       .io_VwirePorts_3_12_5_out( VwireModule_io_VwirePorts_3_12_5_out ),
       .io_VwirePorts_3_12_4_in( ArrayRowModule_3_io_V_wire_out_196 ),
       .io_VwirePorts_3_12_4_en( T1300 ),
       .io_VwirePorts_3_12_4_out( VwireModule_io_VwirePorts_3_12_4_out ),
       .io_VwirePorts_3_12_3_in( ArrayRowModule_3_io_V_wire_out_195 ),
       .io_VwirePorts_3_12_3_en( T1299 ),
       .io_VwirePorts_3_12_3_out( VwireModule_io_VwirePorts_3_12_3_out ),
       .io_VwirePorts_3_12_2_in( ArrayRowModule_3_io_V_wire_out_194 ),
       .io_VwirePorts_3_12_2_en( T1298 ),
       .io_VwirePorts_3_12_2_out( VwireModule_io_VwirePorts_3_12_2_out ),
       .io_VwirePorts_3_12_1_in( ArrayRowModule_3_io_V_wire_out_193 ),
       .io_VwirePorts_3_12_1_en( T1297 ),
       .io_VwirePorts_3_12_1_out( VwireModule_io_VwirePorts_3_12_1_out ),
       .io_VwirePorts_3_12_0_in( ArrayRowModule_3_io_V_wire_out_192 ),
       .io_VwirePorts_3_12_0_en( T1296 ),
       .io_VwirePorts_3_12_0_out( VwireModule_io_VwirePorts_3_12_0_out ),
       .io_VwirePorts_3_11_15_in( ArrayRowModule_3_io_V_wire_out_191 ),
       .io_VwirePorts_3_11_15_en( T1295 ),
       .io_VwirePorts_3_11_15_out( VwireModule_io_VwirePorts_3_11_15_out ),
       .io_VwirePorts_3_11_14_in( ArrayRowModule_3_io_V_wire_out_190 ),
       .io_VwirePorts_3_11_14_en( T1294 ),
       .io_VwirePorts_3_11_14_out( VwireModule_io_VwirePorts_3_11_14_out ),
       .io_VwirePorts_3_11_13_in( ArrayRowModule_3_io_V_wire_out_189 ),
       .io_VwirePorts_3_11_13_en( T1293 ),
       .io_VwirePorts_3_11_13_out( VwireModule_io_VwirePorts_3_11_13_out ),
       .io_VwirePorts_3_11_12_in( ArrayRowModule_3_io_V_wire_out_188 ),
       .io_VwirePorts_3_11_12_en( T1292 ),
       .io_VwirePorts_3_11_12_out( VwireModule_io_VwirePorts_3_11_12_out ),
       .io_VwirePorts_3_11_11_in( ArrayRowModule_3_io_V_wire_out_187 ),
       .io_VwirePorts_3_11_11_en( T1291 ),
       .io_VwirePorts_3_11_11_out( VwireModule_io_VwirePorts_3_11_11_out ),
       .io_VwirePorts_3_11_10_in( ArrayRowModule_3_io_V_wire_out_186 ),
       .io_VwirePorts_3_11_10_en( T1290 ),
       .io_VwirePorts_3_11_10_out( VwireModule_io_VwirePorts_3_11_10_out ),
       .io_VwirePorts_3_11_9_in( ArrayRowModule_3_io_V_wire_out_185 ),
       .io_VwirePorts_3_11_9_en( T1289 ),
       .io_VwirePorts_3_11_9_out( VwireModule_io_VwirePorts_3_11_9_out ),
       .io_VwirePorts_3_11_8_in( ArrayRowModule_3_io_V_wire_out_184 ),
       .io_VwirePorts_3_11_8_en( T1288 ),
       .io_VwirePorts_3_11_8_out( VwireModule_io_VwirePorts_3_11_8_out ),
       .io_VwirePorts_3_11_7_in( ArrayRowModule_3_io_V_wire_out_183 ),
       .io_VwirePorts_3_11_7_en( T1287 ),
       .io_VwirePorts_3_11_7_out( VwireModule_io_VwirePorts_3_11_7_out ),
       .io_VwirePorts_3_11_6_in( ArrayRowModule_3_io_V_wire_out_182 ),
       .io_VwirePorts_3_11_6_en( T1286 ),
       .io_VwirePorts_3_11_6_out( VwireModule_io_VwirePorts_3_11_6_out ),
       .io_VwirePorts_3_11_5_in( ArrayRowModule_3_io_V_wire_out_181 ),
       .io_VwirePorts_3_11_5_en( T1285 ),
       .io_VwirePorts_3_11_5_out( VwireModule_io_VwirePorts_3_11_5_out ),
       .io_VwirePorts_3_11_4_in( ArrayRowModule_3_io_V_wire_out_180 ),
       .io_VwirePorts_3_11_4_en( T1284 ),
       .io_VwirePorts_3_11_4_out( VwireModule_io_VwirePorts_3_11_4_out ),
       .io_VwirePorts_3_11_3_in( ArrayRowModule_3_io_V_wire_out_179 ),
       .io_VwirePorts_3_11_3_en( T1283 ),
       .io_VwirePorts_3_11_3_out( VwireModule_io_VwirePorts_3_11_3_out ),
       .io_VwirePorts_3_11_2_in( ArrayRowModule_3_io_V_wire_out_178 ),
       .io_VwirePorts_3_11_2_en( T1282 ),
       .io_VwirePorts_3_11_2_out( VwireModule_io_VwirePorts_3_11_2_out ),
       .io_VwirePorts_3_11_1_in( ArrayRowModule_3_io_V_wire_out_177 ),
       .io_VwirePorts_3_11_1_en( T1281 ),
       .io_VwirePorts_3_11_1_out( VwireModule_io_VwirePorts_3_11_1_out ),
       .io_VwirePorts_3_11_0_in( ArrayRowModule_3_io_V_wire_out_176 ),
       .io_VwirePorts_3_11_0_en( T1280 ),
       .io_VwirePorts_3_11_0_out( VwireModule_io_VwirePorts_3_11_0_out ),
       .io_VwirePorts_3_10_15_in( ArrayRowModule_3_io_V_wire_out_175 ),
       .io_VwirePorts_3_10_15_en( T1279 ),
       .io_VwirePorts_3_10_15_out( VwireModule_io_VwirePorts_3_10_15_out ),
       .io_VwirePorts_3_10_14_in( ArrayRowModule_3_io_V_wire_out_174 ),
       .io_VwirePorts_3_10_14_en( T1278 ),
       .io_VwirePorts_3_10_14_out( VwireModule_io_VwirePorts_3_10_14_out ),
       .io_VwirePorts_3_10_13_in( ArrayRowModule_3_io_V_wire_out_173 ),
       .io_VwirePorts_3_10_13_en( T1277 ),
       .io_VwirePorts_3_10_13_out( VwireModule_io_VwirePorts_3_10_13_out ),
       .io_VwirePorts_3_10_12_in( ArrayRowModule_3_io_V_wire_out_172 ),
       .io_VwirePorts_3_10_12_en( T1276 ),
       .io_VwirePorts_3_10_12_out( VwireModule_io_VwirePorts_3_10_12_out ),
       .io_VwirePorts_3_10_11_in( ArrayRowModule_3_io_V_wire_out_171 ),
       .io_VwirePorts_3_10_11_en( T1275 ),
       .io_VwirePorts_3_10_11_out( VwireModule_io_VwirePorts_3_10_11_out ),
       .io_VwirePorts_3_10_10_in( ArrayRowModule_3_io_V_wire_out_170 ),
       .io_VwirePorts_3_10_10_en( T1274 ),
       .io_VwirePorts_3_10_10_out( VwireModule_io_VwirePorts_3_10_10_out ),
       .io_VwirePorts_3_10_9_in( ArrayRowModule_3_io_V_wire_out_169 ),
       .io_VwirePorts_3_10_9_en( T1273 ),
       .io_VwirePorts_3_10_9_out( VwireModule_io_VwirePorts_3_10_9_out ),
       .io_VwirePorts_3_10_8_in( ArrayRowModule_3_io_V_wire_out_168 ),
       .io_VwirePorts_3_10_8_en( T1272 ),
       .io_VwirePorts_3_10_8_out( VwireModule_io_VwirePorts_3_10_8_out ),
       .io_VwirePorts_3_10_7_in( ArrayRowModule_3_io_V_wire_out_167 ),
       .io_VwirePorts_3_10_7_en( T1271 ),
       .io_VwirePorts_3_10_7_out( VwireModule_io_VwirePorts_3_10_7_out ),
       .io_VwirePorts_3_10_6_in( ArrayRowModule_3_io_V_wire_out_166 ),
       .io_VwirePorts_3_10_6_en( T1270 ),
       .io_VwirePorts_3_10_6_out( VwireModule_io_VwirePorts_3_10_6_out ),
       .io_VwirePorts_3_10_5_in( ArrayRowModule_3_io_V_wire_out_165 ),
       .io_VwirePorts_3_10_5_en( T1269 ),
       .io_VwirePorts_3_10_5_out( VwireModule_io_VwirePorts_3_10_5_out ),
       .io_VwirePorts_3_10_4_in( ArrayRowModule_3_io_V_wire_out_164 ),
       .io_VwirePorts_3_10_4_en( T1268 ),
       .io_VwirePorts_3_10_4_out( VwireModule_io_VwirePorts_3_10_4_out ),
       .io_VwirePorts_3_10_3_in( ArrayRowModule_3_io_V_wire_out_163 ),
       .io_VwirePorts_3_10_3_en( T1267 ),
       .io_VwirePorts_3_10_3_out( VwireModule_io_VwirePorts_3_10_3_out ),
       .io_VwirePorts_3_10_2_in( ArrayRowModule_3_io_V_wire_out_162 ),
       .io_VwirePorts_3_10_2_en( T1266 ),
       .io_VwirePorts_3_10_2_out( VwireModule_io_VwirePorts_3_10_2_out ),
       .io_VwirePorts_3_10_1_in( ArrayRowModule_3_io_V_wire_out_161 ),
       .io_VwirePorts_3_10_1_en( T1265 ),
       .io_VwirePorts_3_10_1_out( VwireModule_io_VwirePorts_3_10_1_out ),
       .io_VwirePorts_3_10_0_in( ArrayRowModule_3_io_V_wire_out_160 ),
       .io_VwirePorts_3_10_0_en( T1264 ),
       .io_VwirePorts_3_10_0_out( VwireModule_io_VwirePorts_3_10_0_out ),
       .io_VwirePorts_3_9_15_in( ArrayRowModule_3_io_V_wire_out_159 ),
       .io_VwirePorts_3_9_15_en( T1263 ),
       .io_VwirePorts_3_9_15_out( VwireModule_io_VwirePorts_3_9_15_out ),
       .io_VwirePorts_3_9_14_in( ArrayRowModule_3_io_V_wire_out_158 ),
       .io_VwirePorts_3_9_14_en( T1262 ),
       .io_VwirePorts_3_9_14_out( VwireModule_io_VwirePorts_3_9_14_out ),
       .io_VwirePorts_3_9_13_in( ArrayRowModule_3_io_V_wire_out_157 ),
       .io_VwirePorts_3_9_13_en( T1261 ),
       .io_VwirePorts_3_9_13_out( VwireModule_io_VwirePorts_3_9_13_out ),
       .io_VwirePorts_3_9_12_in( ArrayRowModule_3_io_V_wire_out_156 ),
       .io_VwirePorts_3_9_12_en( T1260 ),
       .io_VwirePorts_3_9_12_out( VwireModule_io_VwirePorts_3_9_12_out ),
       .io_VwirePorts_3_9_11_in( ArrayRowModule_3_io_V_wire_out_155 ),
       .io_VwirePorts_3_9_11_en( T1259 ),
       .io_VwirePorts_3_9_11_out( VwireModule_io_VwirePorts_3_9_11_out ),
       .io_VwirePorts_3_9_10_in( ArrayRowModule_3_io_V_wire_out_154 ),
       .io_VwirePorts_3_9_10_en( T1258 ),
       .io_VwirePorts_3_9_10_out( VwireModule_io_VwirePorts_3_9_10_out ),
       .io_VwirePorts_3_9_9_in( ArrayRowModule_3_io_V_wire_out_153 ),
       .io_VwirePorts_3_9_9_en( T1257 ),
       .io_VwirePorts_3_9_9_out( VwireModule_io_VwirePorts_3_9_9_out ),
       .io_VwirePorts_3_9_8_in( ArrayRowModule_3_io_V_wire_out_152 ),
       .io_VwirePorts_3_9_8_en( T1256 ),
       .io_VwirePorts_3_9_8_out( VwireModule_io_VwirePorts_3_9_8_out ),
       .io_VwirePorts_3_9_7_in( ArrayRowModule_3_io_V_wire_out_151 ),
       .io_VwirePorts_3_9_7_en( T1255 ),
       .io_VwirePorts_3_9_7_out( VwireModule_io_VwirePorts_3_9_7_out ),
       .io_VwirePorts_3_9_6_in( ArrayRowModule_3_io_V_wire_out_150 ),
       .io_VwirePorts_3_9_6_en( T1254 ),
       .io_VwirePorts_3_9_6_out( VwireModule_io_VwirePorts_3_9_6_out ),
       .io_VwirePorts_3_9_5_in( ArrayRowModule_3_io_V_wire_out_149 ),
       .io_VwirePorts_3_9_5_en( T1253 ),
       .io_VwirePorts_3_9_5_out( VwireModule_io_VwirePorts_3_9_5_out ),
       .io_VwirePorts_3_9_4_in( ArrayRowModule_3_io_V_wire_out_148 ),
       .io_VwirePorts_3_9_4_en( T1252 ),
       .io_VwirePorts_3_9_4_out( VwireModule_io_VwirePorts_3_9_4_out ),
       .io_VwirePorts_3_9_3_in( ArrayRowModule_3_io_V_wire_out_147 ),
       .io_VwirePorts_3_9_3_en( T1251 ),
       .io_VwirePorts_3_9_3_out( VwireModule_io_VwirePorts_3_9_3_out ),
       .io_VwirePorts_3_9_2_in( ArrayRowModule_3_io_V_wire_out_146 ),
       .io_VwirePorts_3_9_2_en( T1250 ),
       .io_VwirePorts_3_9_2_out( VwireModule_io_VwirePorts_3_9_2_out ),
       .io_VwirePorts_3_9_1_in( ArrayRowModule_3_io_V_wire_out_145 ),
       .io_VwirePorts_3_9_1_en( T1249 ),
       .io_VwirePorts_3_9_1_out( VwireModule_io_VwirePorts_3_9_1_out ),
       .io_VwirePorts_3_9_0_in( ArrayRowModule_3_io_V_wire_out_144 ),
       .io_VwirePorts_3_9_0_en( T1248 ),
       .io_VwirePorts_3_9_0_out( VwireModule_io_VwirePorts_3_9_0_out ),
       .io_VwirePorts_3_8_15_in( ArrayRowModule_3_io_V_wire_out_143 ),
       .io_VwirePorts_3_8_15_en( T1247 ),
       .io_VwirePorts_3_8_15_out( VwireModule_io_VwirePorts_3_8_15_out ),
       .io_VwirePorts_3_8_14_in( ArrayRowModule_3_io_V_wire_out_142 ),
       .io_VwirePorts_3_8_14_en( T1246 ),
       .io_VwirePorts_3_8_14_out( VwireModule_io_VwirePorts_3_8_14_out ),
       .io_VwirePorts_3_8_13_in( ArrayRowModule_3_io_V_wire_out_141 ),
       .io_VwirePorts_3_8_13_en( T1245 ),
       .io_VwirePorts_3_8_13_out( VwireModule_io_VwirePorts_3_8_13_out ),
       .io_VwirePorts_3_8_12_in( ArrayRowModule_3_io_V_wire_out_140 ),
       .io_VwirePorts_3_8_12_en( T1244 ),
       .io_VwirePorts_3_8_12_out( VwireModule_io_VwirePorts_3_8_12_out ),
       .io_VwirePorts_3_8_11_in( ArrayRowModule_3_io_V_wire_out_139 ),
       .io_VwirePorts_3_8_11_en( T1243 ),
       .io_VwirePorts_3_8_11_out( VwireModule_io_VwirePorts_3_8_11_out ),
       .io_VwirePorts_3_8_10_in( ArrayRowModule_3_io_V_wire_out_138 ),
       .io_VwirePorts_3_8_10_en( T1242 ),
       .io_VwirePorts_3_8_10_out( VwireModule_io_VwirePorts_3_8_10_out ),
       .io_VwirePorts_3_8_9_in( ArrayRowModule_3_io_V_wire_out_137 ),
       .io_VwirePorts_3_8_9_en( T1241 ),
       .io_VwirePorts_3_8_9_out( VwireModule_io_VwirePorts_3_8_9_out ),
       .io_VwirePorts_3_8_8_in( ArrayRowModule_3_io_V_wire_out_136 ),
       .io_VwirePorts_3_8_8_en( T1240 ),
       .io_VwirePorts_3_8_8_out( VwireModule_io_VwirePorts_3_8_8_out ),
       .io_VwirePorts_3_8_7_in( ArrayRowModule_3_io_V_wire_out_135 ),
       .io_VwirePorts_3_8_7_en( T1239 ),
       .io_VwirePorts_3_8_7_out( VwireModule_io_VwirePorts_3_8_7_out ),
       .io_VwirePorts_3_8_6_in( ArrayRowModule_3_io_V_wire_out_134 ),
       .io_VwirePorts_3_8_6_en( T1238 ),
       .io_VwirePorts_3_8_6_out( VwireModule_io_VwirePorts_3_8_6_out ),
       .io_VwirePorts_3_8_5_in( ArrayRowModule_3_io_V_wire_out_133 ),
       .io_VwirePorts_3_8_5_en( T1237 ),
       .io_VwirePorts_3_8_5_out( VwireModule_io_VwirePorts_3_8_5_out ),
       .io_VwirePorts_3_8_4_in( ArrayRowModule_3_io_V_wire_out_132 ),
       .io_VwirePorts_3_8_4_en( T1236 ),
       .io_VwirePorts_3_8_4_out( VwireModule_io_VwirePorts_3_8_4_out ),
       .io_VwirePorts_3_8_3_in( ArrayRowModule_3_io_V_wire_out_131 ),
       .io_VwirePorts_3_8_3_en( T1235 ),
       .io_VwirePorts_3_8_3_out( VwireModule_io_VwirePorts_3_8_3_out ),
       .io_VwirePorts_3_8_2_in( ArrayRowModule_3_io_V_wire_out_130 ),
       .io_VwirePorts_3_8_2_en( T1234 ),
       .io_VwirePorts_3_8_2_out( VwireModule_io_VwirePorts_3_8_2_out ),
       .io_VwirePorts_3_8_1_in( ArrayRowModule_3_io_V_wire_out_129 ),
       .io_VwirePorts_3_8_1_en( T1233 ),
       .io_VwirePorts_3_8_1_out( VwireModule_io_VwirePorts_3_8_1_out ),
       .io_VwirePorts_3_8_0_in( ArrayRowModule_3_io_V_wire_out_128 ),
       .io_VwirePorts_3_8_0_en( T1232 ),
       .io_VwirePorts_3_8_0_out( VwireModule_io_VwirePorts_3_8_0_out ),
       .io_VwirePorts_3_7_15_in( ArrayRowModule_3_io_V_wire_out_127 ),
       .io_VwirePorts_3_7_15_en( T1231 ),
       .io_VwirePorts_3_7_15_out( VwireModule_io_VwirePorts_3_7_15_out ),
       .io_VwirePorts_3_7_14_in( ArrayRowModule_3_io_V_wire_out_126 ),
       .io_VwirePorts_3_7_14_en( T1230 ),
       .io_VwirePorts_3_7_14_out( VwireModule_io_VwirePorts_3_7_14_out ),
       .io_VwirePorts_3_7_13_in( ArrayRowModule_3_io_V_wire_out_125 ),
       .io_VwirePorts_3_7_13_en( T1229 ),
       .io_VwirePorts_3_7_13_out( VwireModule_io_VwirePorts_3_7_13_out ),
       .io_VwirePorts_3_7_12_in( ArrayRowModule_3_io_V_wire_out_124 ),
       .io_VwirePorts_3_7_12_en( T1228 ),
       .io_VwirePorts_3_7_12_out( VwireModule_io_VwirePorts_3_7_12_out ),
       .io_VwirePorts_3_7_11_in( ArrayRowModule_3_io_V_wire_out_123 ),
       .io_VwirePorts_3_7_11_en( T1227 ),
       .io_VwirePorts_3_7_11_out( VwireModule_io_VwirePorts_3_7_11_out ),
       .io_VwirePorts_3_7_10_in( ArrayRowModule_3_io_V_wire_out_122 ),
       .io_VwirePorts_3_7_10_en( T1226 ),
       .io_VwirePorts_3_7_10_out( VwireModule_io_VwirePorts_3_7_10_out ),
       .io_VwirePorts_3_7_9_in( ArrayRowModule_3_io_V_wire_out_121 ),
       .io_VwirePorts_3_7_9_en( T1225 ),
       .io_VwirePorts_3_7_9_out( VwireModule_io_VwirePorts_3_7_9_out ),
       .io_VwirePorts_3_7_8_in( ArrayRowModule_3_io_V_wire_out_120 ),
       .io_VwirePorts_3_7_8_en( T1224 ),
       .io_VwirePorts_3_7_8_out( VwireModule_io_VwirePorts_3_7_8_out ),
       .io_VwirePorts_3_7_7_in( ArrayRowModule_3_io_V_wire_out_119 ),
       .io_VwirePorts_3_7_7_en( T1223 ),
       .io_VwirePorts_3_7_7_out( VwireModule_io_VwirePorts_3_7_7_out ),
       .io_VwirePorts_3_7_6_in( ArrayRowModule_3_io_V_wire_out_118 ),
       .io_VwirePorts_3_7_6_en( T1222 ),
       .io_VwirePorts_3_7_6_out( VwireModule_io_VwirePorts_3_7_6_out ),
       .io_VwirePorts_3_7_5_in( ArrayRowModule_3_io_V_wire_out_117 ),
       .io_VwirePorts_3_7_5_en( T1221 ),
       .io_VwirePorts_3_7_5_out( VwireModule_io_VwirePorts_3_7_5_out ),
       .io_VwirePorts_3_7_4_in( ArrayRowModule_3_io_V_wire_out_116 ),
       .io_VwirePorts_3_7_4_en( T1220 ),
       .io_VwirePorts_3_7_4_out( VwireModule_io_VwirePorts_3_7_4_out ),
       .io_VwirePorts_3_7_3_in( ArrayRowModule_3_io_V_wire_out_115 ),
       .io_VwirePorts_3_7_3_en( T1219 ),
       .io_VwirePorts_3_7_3_out( VwireModule_io_VwirePorts_3_7_3_out ),
       .io_VwirePorts_3_7_2_in( ArrayRowModule_3_io_V_wire_out_114 ),
       .io_VwirePorts_3_7_2_en( T1218 ),
       .io_VwirePorts_3_7_2_out( VwireModule_io_VwirePorts_3_7_2_out ),
       .io_VwirePorts_3_7_1_in( ArrayRowModule_3_io_V_wire_out_113 ),
       .io_VwirePorts_3_7_1_en( T1217 ),
       .io_VwirePorts_3_7_1_out( VwireModule_io_VwirePorts_3_7_1_out ),
       .io_VwirePorts_3_7_0_in( ArrayRowModule_3_io_V_wire_out_112 ),
       .io_VwirePorts_3_7_0_en( T1216 ),
       .io_VwirePorts_3_7_0_out( VwireModule_io_VwirePorts_3_7_0_out ),
       .io_VwirePorts_3_6_15_in( ArrayRowModule_3_io_V_wire_out_111 ),
       .io_VwirePorts_3_6_15_en( T1215 ),
       .io_VwirePorts_3_6_15_out( VwireModule_io_VwirePorts_3_6_15_out ),
       .io_VwirePorts_3_6_14_in( ArrayRowModule_3_io_V_wire_out_110 ),
       .io_VwirePorts_3_6_14_en( T1214 ),
       .io_VwirePorts_3_6_14_out( VwireModule_io_VwirePorts_3_6_14_out ),
       .io_VwirePorts_3_6_13_in( ArrayRowModule_3_io_V_wire_out_109 ),
       .io_VwirePorts_3_6_13_en( T1213 ),
       .io_VwirePorts_3_6_13_out( VwireModule_io_VwirePorts_3_6_13_out ),
       .io_VwirePorts_3_6_12_in( ArrayRowModule_3_io_V_wire_out_108 ),
       .io_VwirePorts_3_6_12_en( T1212 ),
       .io_VwirePorts_3_6_12_out( VwireModule_io_VwirePorts_3_6_12_out ),
       .io_VwirePorts_3_6_11_in( ArrayRowModule_3_io_V_wire_out_107 ),
       .io_VwirePorts_3_6_11_en( T1211 ),
       .io_VwirePorts_3_6_11_out( VwireModule_io_VwirePorts_3_6_11_out ),
       .io_VwirePorts_3_6_10_in( ArrayRowModule_3_io_V_wire_out_106 ),
       .io_VwirePorts_3_6_10_en( T1210 ),
       .io_VwirePorts_3_6_10_out( VwireModule_io_VwirePorts_3_6_10_out ),
       .io_VwirePorts_3_6_9_in( ArrayRowModule_3_io_V_wire_out_105 ),
       .io_VwirePorts_3_6_9_en( T1209 ),
       .io_VwirePorts_3_6_9_out( VwireModule_io_VwirePorts_3_6_9_out ),
       .io_VwirePorts_3_6_8_in( ArrayRowModule_3_io_V_wire_out_104 ),
       .io_VwirePorts_3_6_8_en( T1208 ),
       .io_VwirePorts_3_6_8_out( VwireModule_io_VwirePorts_3_6_8_out ),
       .io_VwirePorts_3_6_7_in( ArrayRowModule_3_io_V_wire_out_103 ),
       .io_VwirePorts_3_6_7_en( T1207 ),
       .io_VwirePorts_3_6_7_out( VwireModule_io_VwirePorts_3_6_7_out ),
       .io_VwirePorts_3_6_6_in( ArrayRowModule_3_io_V_wire_out_102 ),
       .io_VwirePorts_3_6_6_en( T1206 ),
       .io_VwirePorts_3_6_6_out( VwireModule_io_VwirePorts_3_6_6_out ),
       .io_VwirePorts_3_6_5_in( ArrayRowModule_3_io_V_wire_out_101 ),
       .io_VwirePorts_3_6_5_en( T1205 ),
       .io_VwirePorts_3_6_5_out( VwireModule_io_VwirePorts_3_6_5_out ),
       .io_VwirePorts_3_6_4_in( ArrayRowModule_3_io_V_wire_out_100 ),
       .io_VwirePorts_3_6_4_en( T1204 ),
       .io_VwirePorts_3_6_4_out( VwireModule_io_VwirePorts_3_6_4_out ),
       .io_VwirePorts_3_6_3_in( ArrayRowModule_3_io_V_wire_out_99 ),
       .io_VwirePorts_3_6_3_en( T1203 ),
       .io_VwirePorts_3_6_3_out( VwireModule_io_VwirePorts_3_6_3_out ),
       .io_VwirePorts_3_6_2_in( ArrayRowModule_3_io_V_wire_out_98 ),
       .io_VwirePorts_3_6_2_en( T1202 ),
       .io_VwirePorts_3_6_2_out( VwireModule_io_VwirePorts_3_6_2_out ),
       .io_VwirePorts_3_6_1_in( ArrayRowModule_3_io_V_wire_out_97 ),
       .io_VwirePorts_3_6_1_en( T1201 ),
       .io_VwirePorts_3_6_1_out( VwireModule_io_VwirePorts_3_6_1_out ),
       .io_VwirePorts_3_6_0_in( ArrayRowModule_3_io_V_wire_out_96 ),
       .io_VwirePorts_3_6_0_en( T1200 ),
       .io_VwirePorts_3_6_0_out( VwireModule_io_VwirePorts_3_6_0_out ),
       .io_VwirePorts_3_5_15_in( ArrayRowModule_3_io_V_wire_out_95 ),
       .io_VwirePorts_3_5_15_en( T1199 ),
       .io_VwirePorts_3_5_15_out( VwireModule_io_VwirePorts_3_5_15_out ),
       .io_VwirePorts_3_5_14_in( ArrayRowModule_3_io_V_wire_out_94 ),
       .io_VwirePorts_3_5_14_en( T1198 ),
       .io_VwirePorts_3_5_14_out( VwireModule_io_VwirePorts_3_5_14_out ),
       .io_VwirePorts_3_5_13_in( ArrayRowModule_3_io_V_wire_out_93 ),
       .io_VwirePorts_3_5_13_en( T1197 ),
       .io_VwirePorts_3_5_13_out( VwireModule_io_VwirePorts_3_5_13_out ),
       .io_VwirePorts_3_5_12_in( ArrayRowModule_3_io_V_wire_out_92 ),
       .io_VwirePorts_3_5_12_en( T1196 ),
       .io_VwirePorts_3_5_12_out( VwireModule_io_VwirePorts_3_5_12_out ),
       .io_VwirePorts_3_5_11_in( ArrayRowModule_3_io_V_wire_out_91 ),
       .io_VwirePorts_3_5_11_en( T1195 ),
       .io_VwirePorts_3_5_11_out( VwireModule_io_VwirePorts_3_5_11_out ),
       .io_VwirePorts_3_5_10_in( ArrayRowModule_3_io_V_wire_out_90 ),
       .io_VwirePorts_3_5_10_en( T1194 ),
       .io_VwirePorts_3_5_10_out( VwireModule_io_VwirePorts_3_5_10_out ),
       .io_VwirePorts_3_5_9_in( ArrayRowModule_3_io_V_wire_out_89 ),
       .io_VwirePorts_3_5_9_en( T1193 ),
       .io_VwirePorts_3_5_9_out( VwireModule_io_VwirePorts_3_5_9_out ),
       .io_VwirePorts_3_5_8_in( ArrayRowModule_3_io_V_wire_out_88 ),
       .io_VwirePorts_3_5_8_en( T1192 ),
       .io_VwirePorts_3_5_8_out( VwireModule_io_VwirePorts_3_5_8_out ),
       .io_VwirePorts_3_5_7_in( ArrayRowModule_3_io_V_wire_out_87 ),
       .io_VwirePorts_3_5_7_en( T1191 ),
       .io_VwirePorts_3_5_7_out( VwireModule_io_VwirePorts_3_5_7_out ),
       .io_VwirePorts_3_5_6_in( ArrayRowModule_3_io_V_wire_out_86 ),
       .io_VwirePorts_3_5_6_en( T1190 ),
       .io_VwirePorts_3_5_6_out( VwireModule_io_VwirePorts_3_5_6_out ),
       .io_VwirePorts_3_5_5_in( ArrayRowModule_3_io_V_wire_out_85 ),
       .io_VwirePorts_3_5_5_en( T1189 ),
       .io_VwirePorts_3_5_5_out( VwireModule_io_VwirePorts_3_5_5_out ),
       .io_VwirePorts_3_5_4_in( ArrayRowModule_3_io_V_wire_out_84 ),
       .io_VwirePorts_3_5_4_en( T1188 ),
       .io_VwirePorts_3_5_4_out( VwireModule_io_VwirePorts_3_5_4_out ),
       .io_VwirePorts_3_5_3_in( ArrayRowModule_3_io_V_wire_out_83 ),
       .io_VwirePorts_3_5_3_en( T1187 ),
       .io_VwirePorts_3_5_3_out( VwireModule_io_VwirePorts_3_5_3_out ),
       .io_VwirePorts_3_5_2_in( ArrayRowModule_3_io_V_wire_out_82 ),
       .io_VwirePorts_3_5_2_en( T1186 ),
       .io_VwirePorts_3_5_2_out( VwireModule_io_VwirePorts_3_5_2_out ),
       .io_VwirePorts_3_5_1_in( ArrayRowModule_3_io_V_wire_out_81 ),
       .io_VwirePorts_3_5_1_en( T1185 ),
       .io_VwirePorts_3_5_1_out( VwireModule_io_VwirePorts_3_5_1_out ),
       .io_VwirePorts_3_5_0_in( ArrayRowModule_3_io_V_wire_out_80 ),
       .io_VwirePorts_3_5_0_en( T1184 ),
       .io_VwirePorts_3_5_0_out( VwireModule_io_VwirePorts_3_5_0_out ),
       .io_VwirePorts_3_4_15_in( ArrayRowModule_3_io_V_wire_out_79 ),
       .io_VwirePorts_3_4_15_en( T1183 ),
       .io_VwirePorts_3_4_15_out( VwireModule_io_VwirePorts_3_4_15_out ),
       .io_VwirePorts_3_4_14_in( ArrayRowModule_3_io_V_wire_out_78 ),
       .io_VwirePorts_3_4_14_en( T1182 ),
       .io_VwirePorts_3_4_14_out( VwireModule_io_VwirePorts_3_4_14_out ),
       .io_VwirePorts_3_4_13_in( ArrayRowModule_3_io_V_wire_out_77 ),
       .io_VwirePorts_3_4_13_en( T1181 ),
       .io_VwirePorts_3_4_13_out( VwireModule_io_VwirePorts_3_4_13_out ),
       .io_VwirePorts_3_4_12_in( ArrayRowModule_3_io_V_wire_out_76 ),
       .io_VwirePorts_3_4_12_en( T1180 ),
       .io_VwirePorts_3_4_12_out( VwireModule_io_VwirePorts_3_4_12_out ),
       .io_VwirePorts_3_4_11_in( ArrayRowModule_3_io_V_wire_out_75 ),
       .io_VwirePorts_3_4_11_en( T1179 ),
       .io_VwirePorts_3_4_11_out( VwireModule_io_VwirePorts_3_4_11_out ),
       .io_VwirePorts_3_4_10_in( ArrayRowModule_3_io_V_wire_out_74 ),
       .io_VwirePorts_3_4_10_en( T1178 ),
       .io_VwirePorts_3_4_10_out( VwireModule_io_VwirePorts_3_4_10_out ),
       .io_VwirePorts_3_4_9_in( ArrayRowModule_3_io_V_wire_out_73 ),
       .io_VwirePorts_3_4_9_en( T1177 ),
       .io_VwirePorts_3_4_9_out( VwireModule_io_VwirePorts_3_4_9_out ),
       .io_VwirePorts_3_4_8_in( ArrayRowModule_3_io_V_wire_out_72 ),
       .io_VwirePorts_3_4_8_en( T1176 ),
       .io_VwirePorts_3_4_8_out( VwireModule_io_VwirePorts_3_4_8_out ),
       .io_VwirePorts_3_4_7_in( ArrayRowModule_3_io_V_wire_out_71 ),
       .io_VwirePorts_3_4_7_en( T1175 ),
       .io_VwirePorts_3_4_7_out( VwireModule_io_VwirePorts_3_4_7_out ),
       .io_VwirePorts_3_4_6_in( ArrayRowModule_3_io_V_wire_out_70 ),
       .io_VwirePorts_3_4_6_en( T1174 ),
       .io_VwirePorts_3_4_6_out( VwireModule_io_VwirePorts_3_4_6_out ),
       .io_VwirePorts_3_4_5_in( ArrayRowModule_3_io_V_wire_out_69 ),
       .io_VwirePorts_3_4_5_en( T1173 ),
       .io_VwirePorts_3_4_5_out( VwireModule_io_VwirePorts_3_4_5_out ),
       .io_VwirePorts_3_4_4_in( ArrayRowModule_3_io_V_wire_out_68 ),
       .io_VwirePorts_3_4_4_en( T1172 ),
       .io_VwirePorts_3_4_4_out( VwireModule_io_VwirePorts_3_4_4_out ),
       .io_VwirePorts_3_4_3_in( ArrayRowModule_3_io_V_wire_out_67 ),
       .io_VwirePorts_3_4_3_en( T1171 ),
       .io_VwirePorts_3_4_3_out( VwireModule_io_VwirePorts_3_4_3_out ),
       .io_VwirePorts_3_4_2_in( ArrayRowModule_3_io_V_wire_out_66 ),
       .io_VwirePorts_3_4_2_en( T1170 ),
       .io_VwirePorts_3_4_2_out( VwireModule_io_VwirePorts_3_4_2_out ),
       .io_VwirePorts_3_4_1_in( ArrayRowModule_3_io_V_wire_out_65 ),
       .io_VwirePorts_3_4_1_en( T1169 ),
       .io_VwirePorts_3_4_1_out( VwireModule_io_VwirePorts_3_4_1_out ),
       .io_VwirePorts_3_4_0_in( ArrayRowModule_3_io_V_wire_out_64 ),
       .io_VwirePorts_3_4_0_en( T1168 ),
       .io_VwirePorts_3_4_0_out( VwireModule_io_VwirePorts_3_4_0_out ),
       .io_VwirePorts_3_3_15_in( ArrayRowModule_3_io_V_wire_out_63 ),
       .io_VwirePorts_3_3_15_en( T1167 ),
       .io_VwirePorts_3_3_15_out( VwireModule_io_VwirePorts_3_3_15_out ),
       .io_VwirePorts_3_3_14_in( ArrayRowModule_3_io_V_wire_out_62 ),
       .io_VwirePorts_3_3_14_en( T1166 ),
       .io_VwirePorts_3_3_14_out( VwireModule_io_VwirePorts_3_3_14_out ),
       .io_VwirePorts_3_3_13_in( ArrayRowModule_3_io_V_wire_out_61 ),
       .io_VwirePorts_3_3_13_en( T1165 ),
       .io_VwirePorts_3_3_13_out( VwireModule_io_VwirePorts_3_3_13_out ),
       .io_VwirePorts_3_3_12_in( ArrayRowModule_3_io_V_wire_out_60 ),
       .io_VwirePorts_3_3_12_en( T1164 ),
       .io_VwirePorts_3_3_12_out( VwireModule_io_VwirePorts_3_3_12_out ),
       .io_VwirePorts_3_3_11_in( ArrayRowModule_3_io_V_wire_out_59 ),
       .io_VwirePorts_3_3_11_en( T1163 ),
       .io_VwirePorts_3_3_11_out( VwireModule_io_VwirePorts_3_3_11_out ),
       .io_VwirePorts_3_3_10_in( ArrayRowModule_3_io_V_wire_out_58 ),
       .io_VwirePorts_3_3_10_en( T1162 ),
       .io_VwirePorts_3_3_10_out( VwireModule_io_VwirePorts_3_3_10_out ),
       .io_VwirePorts_3_3_9_in( ArrayRowModule_3_io_V_wire_out_57 ),
       .io_VwirePorts_3_3_9_en( T1161 ),
       .io_VwirePorts_3_3_9_out( VwireModule_io_VwirePorts_3_3_9_out ),
       .io_VwirePorts_3_3_8_in( ArrayRowModule_3_io_V_wire_out_56 ),
       .io_VwirePorts_3_3_8_en( T1160 ),
       .io_VwirePorts_3_3_8_out( VwireModule_io_VwirePorts_3_3_8_out ),
       .io_VwirePorts_3_3_7_in( ArrayRowModule_3_io_V_wire_out_55 ),
       .io_VwirePorts_3_3_7_en( T1159 ),
       .io_VwirePorts_3_3_7_out( VwireModule_io_VwirePorts_3_3_7_out ),
       .io_VwirePorts_3_3_6_in( ArrayRowModule_3_io_V_wire_out_54 ),
       .io_VwirePorts_3_3_6_en( T1158 ),
       .io_VwirePorts_3_3_6_out( VwireModule_io_VwirePorts_3_3_6_out ),
       .io_VwirePorts_3_3_5_in( ArrayRowModule_3_io_V_wire_out_53 ),
       .io_VwirePorts_3_3_5_en( T1157 ),
       .io_VwirePorts_3_3_5_out( VwireModule_io_VwirePorts_3_3_5_out ),
       .io_VwirePorts_3_3_4_in( ArrayRowModule_3_io_V_wire_out_52 ),
       .io_VwirePorts_3_3_4_en( T1156 ),
       .io_VwirePorts_3_3_4_out( VwireModule_io_VwirePorts_3_3_4_out ),
       .io_VwirePorts_3_3_3_in( ArrayRowModule_3_io_V_wire_out_51 ),
       .io_VwirePorts_3_3_3_en( T1155 ),
       .io_VwirePorts_3_3_3_out( VwireModule_io_VwirePorts_3_3_3_out ),
       .io_VwirePorts_3_3_2_in( ArrayRowModule_3_io_V_wire_out_50 ),
       .io_VwirePorts_3_3_2_en( T1154 ),
       .io_VwirePorts_3_3_2_out( VwireModule_io_VwirePorts_3_3_2_out ),
       .io_VwirePorts_3_3_1_in( ArrayRowModule_3_io_V_wire_out_49 ),
       .io_VwirePorts_3_3_1_en( T1153 ),
       .io_VwirePorts_3_3_1_out( VwireModule_io_VwirePorts_3_3_1_out ),
       .io_VwirePorts_3_3_0_in( ArrayRowModule_3_io_V_wire_out_48 ),
       .io_VwirePorts_3_3_0_en( T1152 ),
       .io_VwirePorts_3_3_0_out( VwireModule_io_VwirePorts_3_3_0_out ),
       .io_VwirePorts_3_2_15_in( ArrayRowModule_3_io_V_wire_out_47 ),
       .io_VwirePorts_3_2_15_en( T1151 ),
       .io_VwirePorts_3_2_15_out( VwireModule_io_VwirePorts_3_2_15_out ),
       .io_VwirePorts_3_2_14_in( ArrayRowModule_3_io_V_wire_out_46 ),
       .io_VwirePorts_3_2_14_en( T1150 ),
       .io_VwirePorts_3_2_14_out( VwireModule_io_VwirePorts_3_2_14_out ),
       .io_VwirePorts_3_2_13_in( ArrayRowModule_3_io_V_wire_out_45 ),
       .io_VwirePorts_3_2_13_en( T1149 ),
       .io_VwirePorts_3_2_13_out( VwireModule_io_VwirePorts_3_2_13_out ),
       .io_VwirePorts_3_2_12_in( ArrayRowModule_3_io_V_wire_out_44 ),
       .io_VwirePorts_3_2_12_en( T1148 ),
       .io_VwirePorts_3_2_12_out( VwireModule_io_VwirePorts_3_2_12_out ),
       .io_VwirePorts_3_2_11_in( ArrayRowModule_3_io_V_wire_out_43 ),
       .io_VwirePorts_3_2_11_en( T1147 ),
       .io_VwirePorts_3_2_11_out( VwireModule_io_VwirePorts_3_2_11_out ),
       .io_VwirePorts_3_2_10_in( ArrayRowModule_3_io_V_wire_out_42 ),
       .io_VwirePorts_3_2_10_en( T1146 ),
       .io_VwirePorts_3_2_10_out( VwireModule_io_VwirePorts_3_2_10_out ),
       .io_VwirePorts_3_2_9_in( ArrayRowModule_3_io_V_wire_out_41 ),
       .io_VwirePorts_3_2_9_en( T1145 ),
       .io_VwirePorts_3_2_9_out( VwireModule_io_VwirePorts_3_2_9_out ),
       .io_VwirePorts_3_2_8_in( ArrayRowModule_3_io_V_wire_out_40 ),
       .io_VwirePorts_3_2_8_en( T1144 ),
       .io_VwirePorts_3_2_8_out( VwireModule_io_VwirePorts_3_2_8_out ),
       .io_VwirePorts_3_2_7_in( ArrayRowModule_3_io_V_wire_out_39 ),
       .io_VwirePorts_3_2_7_en( T1143 ),
       .io_VwirePorts_3_2_7_out( VwireModule_io_VwirePorts_3_2_7_out ),
       .io_VwirePorts_3_2_6_in( ArrayRowModule_3_io_V_wire_out_38 ),
       .io_VwirePorts_3_2_6_en( T1142 ),
       .io_VwirePorts_3_2_6_out( VwireModule_io_VwirePorts_3_2_6_out ),
       .io_VwirePorts_3_2_5_in( ArrayRowModule_3_io_V_wire_out_37 ),
       .io_VwirePorts_3_2_5_en( T1141 ),
       .io_VwirePorts_3_2_5_out( VwireModule_io_VwirePorts_3_2_5_out ),
       .io_VwirePorts_3_2_4_in( ArrayRowModule_3_io_V_wire_out_36 ),
       .io_VwirePorts_3_2_4_en( T1140 ),
       .io_VwirePorts_3_2_4_out( VwireModule_io_VwirePorts_3_2_4_out ),
       .io_VwirePorts_3_2_3_in( ArrayRowModule_3_io_V_wire_out_35 ),
       .io_VwirePorts_3_2_3_en( T1139 ),
       .io_VwirePorts_3_2_3_out( VwireModule_io_VwirePorts_3_2_3_out ),
       .io_VwirePorts_3_2_2_in( ArrayRowModule_3_io_V_wire_out_34 ),
       .io_VwirePorts_3_2_2_en( T1138 ),
       .io_VwirePorts_3_2_2_out( VwireModule_io_VwirePorts_3_2_2_out ),
       .io_VwirePorts_3_2_1_in( ArrayRowModule_3_io_V_wire_out_33 ),
       .io_VwirePorts_3_2_1_en( T1137 ),
       .io_VwirePorts_3_2_1_out( VwireModule_io_VwirePorts_3_2_1_out ),
       .io_VwirePorts_3_2_0_in( ArrayRowModule_3_io_V_wire_out_32 ),
       .io_VwirePorts_3_2_0_en( T1136 ),
       .io_VwirePorts_3_2_0_out( VwireModule_io_VwirePorts_3_2_0_out ),
       .io_VwirePorts_3_1_15_in( ArrayRowModule_3_io_V_wire_out_31 ),
       .io_VwirePorts_3_1_15_en( T1135 ),
       .io_VwirePorts_3_1_15_out( VwireModule_io_VwirePorts_3_1_15_out ),
       .io_VwirePorts_3_1_14_in( ArrayRowModule_3_io_V_wire_out_30 ),
       .io_VwirePorts_3_1_14_en( T1134 ),
       .io_VwirePorts_3_1_14_out( VwireModule_io_VwirePorts_3_1_14_out ),
       .io_VwirePorts_3_1_13_in( ArrayRowModule_3_io_V_wire_out_29 ),
       .io_VwirePorts_3_1_13_en( T1133 ),
       .io_VwirePorts_3_1_13_out( VwireModule_io_VwirePorts_3_1_13_out ),
       .io_VwirePorts_3_1_12_in( ArrayRowModule_3_io_V_wire_out_28 ),
       .io_VwirePorts_3_1_12_en( T1132 ),
       .io_VwirePorts_3_1_12_out( VwireModule_io_VwirePorts_3_1_12_out ),
       .io_VwirePorts_3_1_11_in( ArrayRowModule_3_io_V_wire_out_27 ),
       .io_VwirePorts_3_1_11_en( T1131 ),
       .io_VwirePorts_3_1_11_out( VwireModule_io_VwirePorts_3_1_11_out ),
       .io_VwirePorts_3_1_10_in( ArrayRowModule_3_io_V_wire_out_26 ),
       .io_VwirePorts_3_1_10_en( T1130 ),
       .io_VwirePorts_3_1_10_out( VwireModule_io_VwirePorts_3_1_10_out ),
       .io_VwirePorts_3_1_9_in( ArrayRowModule_3_io_V_wire_out_25 ),
       .io_VwirePorts_3_1_9_en( T1129 ),
       .io_VwirePorts_3_1_9_out( VwireModule_io_VwirePorts_3_1_9_out ),
       .io_VwirePorts_3_1_8_in( ArrayRowModule_3_io_V_wire_out_24 ),
       .io_VwirePorts_3_1_8_en( T1128 ),
       .io_VwirePorts_3_1_8_out( VwireModule_io_VwirePorts_3_1_8_out ),
       .io_VwirePorts_3_1_7_in( ArrayRowModule_3_io_V_wire_out_23 ),
       .io_VwirePorts_3_1_7_en( T1127 ),
       .io_VwirePorts_3_1_7_out( VwireModule_io_VwirePorts_3_1_7_out ),
       .io_VwirePorts_3_1_6_in( ArrayRowModule_3_io_V_wire_out_22 ),
       .io_VwirePorts_3_1_6_en( T1126 ),
       .io_VwirePorts_3_1_6_out( VwireModule_io_VwirePorts_3_1_6_out ),
       .io_VwirePorts_3_1_5_in( ArrayRowModule_3_io_V_wire_out_21 ),
       .io_VwirePorts_3_1_5_en( T1125 ),
       .io_VwirePorts_3_1_5_out( VwireModule_io_VwirePorts_3_1_5_out ),
       .io_VwirePorts_3_1_4_in( ArrayRowModule_3_io_V_wire_out_20 ),
       .io_VwirePorts_3_1_4_en( T1124 ),
       .io_VwirePorts_3_1_4_out( VwireModule_io_VwirePorts_3_1_4_out ),
       .io_VwirePorts_3_1_3_in( ArrayRowModule_3_io_V_wire_out_19 ),
       .io_VwirePorts_3_1_3_en( T1123 ),
       .io_VwirePorts_3_1_3_out( VwireModule_io_VwirePorts_3_1_3_out ),
       .io_VwirePorts_3_1_2_in( ArrayRowModule_3_io_V_wire_out_18 ),
       .io_VwirePorts_3_1_2_en( T1122 ),
       .io_VwirePorts_3_1_2_out( VwireModule_io_VwirePorts_3_1_2_out ),
       .io_VwirePorts_3_1_1_in( ArrayRowModule_3_io_V_wire_out_17 ),
       .io_VwirePorts_3_1_1_en( T1121 ),
       .io_VwirePorts_3_1_1_out( VwireModule_io_VwirePorts_3_1_1_out ),
       .io_VwirePorts_3_1_0_in( ArrayRowModule_3_io_V_wire_out_16 ),
       .io_VwirePorts_3_1_0_en( T1120 ),
       .io_VwirePorts_3_1_0_out( VwireModule_io_VwirePorts_3_1_0_out ),
       .io_VwirePorts_3_0_15_in( ArrayRowModule_3_io_V_wire_out_15 ),
       .io_VwirePorts_3_0_15_en( T1119 ),
       .io_VwirePorts_3_0_15_out( VwireModule_io_VwirePorts_3_0_15_out ),
       .io_VwirePorts_3_0_14_in( ArrayRowModule_3_io_V_wire_out_14 ),
       .io_VwirePorts_3_0_14_en( T1118 ),
       .io_VwirePorts_3_0_14_out( VwireModule_io_VwirePorts_3_0_14_out ),
       .io_VwirePorts_3_0_13_in( ArrayRowModule_3_io_V_wire_out_13 ),
       .io_VwirePorts_3_0_13_en( T1117 ),
       .io_VwirePorts_3_0_13_out( VwireModule_io_VwirePorts_3_0_13_out ),
       .io_VwirePorts_3_0_12_in( ArrayRowModule_3_io_V_wire_out_12 ),
       .io_VwirePorts_3_0_12_en( T1116 ),
       .io_VwirePorts_3_0_12_out( VwireModule_io_VwirePorts_3_0_12_out ),
       .io_VwirePorts_3_0_11_in( ArrayRowModule_3_io_V_wire_out_11 ),
       .io_VwirePorts_3_0_11_en( T1115 ),
       .io_VwirePorts_3_0_11_out( VwireModule_io_VwirePorts_3_0_11_out ),
       .io_VwirePorts_3_0_10_in( ArrayRowModule_3_io_V_wire_out_10 ),
       .io_VwirePorts_3_0_10_en( T1114 ),
       .io_VwirePorts_3_0_10_out( VwireModule_io_VwirePorts_3_0_10_out ),
       .io_VwirePorts_3_0_9_in( ArrayRowModule_3_io_V_wire_out_9 ),
       .io_VwirePorts_3_0_9_en( T1113 ),
       .io_VwirePorts_3_0_9_out( VwireModule_io_VwirePorts_3_0_9_out ),
       .io_VwirePorts_3_0_8_in( ArrayRowModule_3_io_V_wire_out_8 ),
       .io_VwirePorts_3_0_8_en( T1112 ),
       .io_VwirePorts_3_0_8_out( VwireModule_io_VwirePorts_3_0_8_out ),
       .io_VwirePorts_3_0_7_in( ArrayRowModule_3_io_V_wire_out_7 ),
       .io_VwirePorts_3_0_7_en( T1111 ),
       .io_VwirePorts_3_0_7_out( VwireModule_io_VwirePorts_3_0_7_out ),
       .io_VwirePorts_3_0_6_in( ArrayRowModule_3_io_V_wire_out_6 ),
       .io_VwirePorts_3_0_6_en( T1110 ),
       .io_VwirePorts_3_0_6_out( VwireModule_io_VwirePorts_3_0_6_out ),
       .io_VwirePorts_3_0_5_in( ArrayRowModule_3_io_V_wire_out_5 ),
       .io_VwirePorts_3_0_5_en( T1109 ),
       .io_VwirePorts_3_0_5_out( VwireModule_io_VwirePorts_3_0_5_out ),
       .io_VwirePorts_3_0_4_in( ArrayRowModule_3_io_V_wire_out_4 ),
       .io_VwirePorts_3_0_4_en( T1108 ),
       .io_VwirePorts_3_0_4_out( VwireModule_io_VwirePorts_3_0_4_out ),
       .io_VwirePorts_3_0_3_in( ArrayRowModule_3_io_V_wire_out_3 ),
       .io_VwirePorts_3_0_3_en( T1107 ),
       .io_VwirePorts_3_0_3_out( VwireModule_io_VwirePorts_3_0_3_out ),
       .io_VwirePorts_3_0_2_in( ArrayRowModule_3_io_V_wire_out_2 ),
       .io_VwirePorts_3_0_2_en( T1106 ),
       .io_VwirePorts_3_0_2_out( VwireModule_io_VwirePorts_3_0_2_out ),
       .io_VwirePorts_3_0_1_in( ArrayRowModule_3_io_V_wire_out_1 ),
       .io_VwirePorts_3_0_1_en( T1105 ),
       .io_VwirePorts_3_0_1_out( VwireModule_io_VwirePorts_3_0_1_out ),
       .io_VwirePorts_3_0_0_in( ArrayRowModule_3_io_V_wire_out_0 ),
       .io_VwirePorts_3_0_0_en( T1104 ),
       .io_VwirePorts_3_0_0_out( VwireModule_io_VwirePorts_3_0_0_out ),
       .io_VwirePorts_2_22_15_in( ArrayRowModule_2_io_V_wire_out_367 ),
       .io_VwirePorts_2_22_15_en( T1103 ),
       .io_VwirePorts_2_22_15_out( VwireModule_io_VwirePorts_2_22_15_out ),
       .io_VwirePorts_2_22_14_in( ArrayRowModule_2_io_V_wire_out_366 ),
       .io_VwirePorts_2_22_14_en( T1102 ),
       .io_VwirePorts_2_22_14_out( VwireModule_io_VwirePorts_2_22_14_out ),
       .io_VwirePorts_2_22_13_in( ArrayRowModule_2_io_V_wire_out_365 ),
       .io_VwirePorts_2_22_13_en( T1101 ),
       .io_VwirePorts_2_22_13_out( VwireModule_io_VwirePorts_2_22_13_out ),
       .io_VwirePorts_2_22_12_in( ArrayRowModule_2_io_V_wire_out_364 ),
       .io_VwirePorts_2_22_12_en( T1100 ),
       .io_VwirePorts_2_22_12_out( VwireModule_io_VwirePorts_2_22_12_out ),
       .io_VwirePorts_2_22_11_in( ArrayRowModule_2_io_V_wire_out_363 ),
       .io_VwirePorts_2_22_11_en( T1099 ),
       .io_VwirePorts_2_22_11_out( VwireModule_io_VwirePorts_2_22_11_out ),
       .io_VwirePorts_2_22_10_in( ArrayRowModule_2_io_V_wire_out_362 ),
       .io_VwirePorts_2_22_10_en( T1098 ),
       .io_VwirePorts_2_22_10_out( VwireModule_io_VwirePorts_2_22_10_out ),
       .io_VwirePorts_2_22_9_in( ArrayRowModule_2_io_V_wire_out_361 ),
       .io_VwirePorts_2_22_9_en( T1097 ),
       .io_VwirePorts_2_22_9_out( VwireModule_io_VwirePorts_2_22_9_out ),
       .io_VwirePorts_2_22_8_in( ArrayRowModule_2_io_V_wire_out_360 ),
       .io_VwirePorts_2_22_8_en( T1096 ),
       .io_VwirePorts_2_22_8_out( VwireModule_io_VwirePorts_2_22_8_out ),
       .io_VwirePorts_2_22_7_in( ArrayRowModule_2_io_V_wire_out_359 ),
       .io_VwirePorts_2_22_7_en( T1095 ),
       .io_VwirePorts_2_22_7_out( VwireModule_io_VwirePorts_2_22_7_out ),
       .io_VwirePorts_2_22_6_in( ArrayRowModule_2_io_V_wire_out_358 ),
       .io_VwirePorts_2_22_6_en( T1094 ),
       .io_VwirePorts_2_22_6_out( VwireModule_io_VwirePorts_2_22_6_out ),
       .io_VwirePorts_2_22_5_in( ArrayRowModule_2_io_V_wire_out_357 ),
       .io_VwirePorts_2_22_5_en( T1093 ),
       .io_VwirePorts_2_22_5_out( VwireModule_io_VwirePorts_2_22_5_out ),
       .io_VwirePorts_2_22_4_in( ArrayRowModule_2_io_V_wire_out_356 ),
       .io_VwirePorts_2_22_4_en( T1092 ),
       .io_VwirePorts_2_22_4_out( VwireModule_io_VwirePorts_2_22_4_out ),
       .io_VwirePorts_2_22_3_in( ArrayRowModule_2_io_V_wire_out_355 ),
       .io_VwirePorts_2_22_3_en( T1091 ),
       .io_VwirePorts_2_22_3_out( VwireModule_io_VwirePorts_2_22_3_out ),
       .io_VwirePorts_2_22_2_in( ArrayRowModule_2_io_V_wire_out_354 ),
       .io_VwirePorts_2_22_2_en( T1090 ),
       .io_VwirePorts_2_22_2_out( VwireModule_io_VwirePorts_2_22_2_out ),
       .io_VwirePorts_2_22_1_in( ArrayRowModule_2_io_V_wire_out_353 ),
       .io_VwirePorts_2_22_1_en( T1089 ),
       .io_VwirePorts_2_22_1_out( VwireModule_io_VwirePorts_2_22_1_out ),
       .io_VwirePorts_2_22_0_in( ArrayRowModule_2_io_V_wire_out_352 ),
       .io_VwirePorts_2_22_0_en( T1088 ),
       .io_VwirePorts_2_22_0_out( VwireModule_io_VwirePorts_2_22_0_out ),
       .io_VwirePorts_2_21_15_in( ArrayRowModule_2_io_V_wire_out_351 ),
       .io_VwirePorts_2_21_15_en( T1087 ),
       .io_VwirePorts_2_21_15_out( VwireModule_io_VwirePorts_2_21_15_out ),
       .io_VwirePorts_2_21_14_in( ArrayRowModule_2_io_V_wire_out_350 ),
       .io_VwirePorts_2_21_14_en( T1086 ),
       .io_VwirePorts_2_21_14_out( VwireModule_io_VwirePorts_2_21_14_out ),
       .io_VwirePorts_2_21_13_in( ArrayRowModule_2_io_V_wire_out_349 ),
       .io_VwirePorts_2_21_13_en( T1085 ),
       .io_VwirePorts_2_21_13_out( VwireModule_io_VwirePorts_2_21_13_out ),
       .io_VwirePorts_2_21_12_in( ArrayRowModule_2_io_V_wire_out_348 ),
       .io_VwirePorts_2_21_12_en( T1084 ),
       .io_VwirePorts_2_21_12_out( VwireModule_io_VwirePorts_2_21_12_out ),
       .io_VwirePorts_2_21_11_in( ArrayRowModule_2_io_V_wire_out_347 ),
       .io_VwirePorts_2_21_11_en( T1083 ),
       .io_VwirePorts_2_21_11_out( VwireModule_io_VwirePorts_2_21_11_out ),
       .io_VwirePorts_2_21_10_in( ArrayRowModule_2_io_V_wire_out_346 ),
       .io_VwirePorts_2_21_10_en( T1082 ),
       .io_VwirePorts_2_21_10_out( VwireModule_io_VwirePorts_2_21_10_out ),
       .io_VwirePorts_2_21_9_in( ArrayRowModule_2_io_V_wire_out_345 ),
       .io_VwirePorts_2_21_9_en( T1081 ),
       .io_VwirePorts_2_21_9_out( VwireModule_io_VwirePorts_2_21_9_out ),
       .io_VwirePorts_2_21_8_in( ArrayRowModule_2_io_V_wire_out_344 ),
       .io_VwirePorts_2_21_8_en( T1080 ),
       .io_VwirePorts_2_21_8_out( VwireModule_io_VwirePorts_2_21_8_out ),
       .io_VwirePorts_2_21_7_in( ArrayRowModule_2_io_V_wire_out_343 ),
       .io_VwirePorts_2_21_7_en( T1079 ),
       .io_VwirePorts_2_21_7_out( VwireModule_io_VwirePorts_2_21_7_out ),
       .io_VwirePorts_2_21_6_in( ArrayRowModule_2_io_V_wire_out_342 ),
       .io_VwirePorts_2_21_6_en( T1078 ),
       .io_VwirePorts_2_21_6_out( VwireModule_io_VwirePorts_2_21_6_out ),
       .io_VwirePorts_2_21_5_in( ArrayRowModule_2_io_V_wire_out_341 ),
       .io_VwirePorts_2_21_5_en( T1077 ),
       .io_VwirePorts_2_21_5_out( VwireModule_io_VwirePorts_2_21_5_out ),
       .io_VwirePorts_2_21_4_in( ArrayRowModule_2_io_V_wire_out_340 ),
       .io_VwirePorts_2_21_4_en( T1076 ),
       .io_VwirePorts_2_21_4_out( VwireModule_io_VwirePorts_2_21_4_out ),
       .io_VwirePorts_2_21_3_in( ArrayRowModule_2_io_V_wire_out_339 ),
       .io_VwirePorts_2_21_3_en( T1075 ),
       .io_VwirePorts_2_21_3_out( VwireModule_io_VwirePorts_2_21_3_out ),
       .io_VwirePorts_2_21_2_in( ArrayRowModule_2_io_V_wire_out_338 ),
       .io_VwirePorts_2_21_2_en( T1074 ),
       .io_VwirePorts_2_21_2_out( VwireModule_io_VwirePorts_2_21_2_out ),
       .io_VwirePorts_2_21_1_in( ArrayRowModule_2_io_V_wire_out_337 ),
       .io_VwirePorts_2_21_1_en( T1073 ),
       .io_VwirePorts_2_21_1_out( VwireModule_io_VwirePorts_2_21_1_out ),
       .io_VwirePorts_2_21_0_in( ArrayRowModule_2_io_V_wire_out_336 ),
       .io_VwirePorts_2_21_0_en( T1072 ),
       .io_VwirePorts_2_21_0_out( VwireModule_io_VwirePorts_2_21_0_out ),
       .io_VwirePorts_2_20_15_in( ArrayRowModule_2_io_V_wire_out_335 ),
       .io_VwirePorts_2_20_15_en( T1071 ),
       .io_VwirePorts_2_20_15_out( VwireModule_io_VwirePorts_2_20_15_out ),
       .io_VwirePorts_2_20_14_in( ArrayRowModule_2_io_V_wire_out_334 ),
       .io_VwirePorts_2_20_14_en( T1070 ),
       .io_VwirePorts_2_20_14_out( VwireModule_io_VwirePorts_2_20_14_out ),
       .io_VwirePorts_2_20_13_in( ArrayRowModule_2_io_V_wire_out_333 ),
       .io_VwirePorts_2_20_13_en( T1069 ),
       .io_VwirePorts_2_20_13_out( VwireModule_io_VwirePorts_2_20_13_out ),
       .io_VwirePorts_2_20_12_in( ArrayRowModule_2_io_V_wire_out_332 ),
       .io_VwirePorts_2_20_12_en( T1068 ),
       .io_VwirePorts_2_20_12_out( VwireModule_io_VwirePorts_2_20_12_out ),
       .io_VwirePorts_2_20_11_in( ArrayRowModule_2_io_V_wire_out_331 ),
       .io_VwirePorts_2_20_11_en( T1067 ),
       .io_VwirePorts_2_20_11_out( VwireModule_io_VwirePorts_2_20_11_out ),
       .io_VwirePorts_2_20_10_in( ArrayRowModule_2_io_V_wire_out_330 ),
       .io_VwirePorts_2_20_10_en( T1066 ),
       .io_VwirePorts_2_20_10_out( VwireModule_io_VwirePorts_2_20_10_out ),
       .io_VwirePorts_2_20_9_in( ArrayRowModule_2_io_V_wire_out_329 ),
       .io_VwirePorts_2_20_9_en( T1065 ),
       .io_VwirePorts_2_20_9_out( VwireModule_io_VwirePorts_2_20_9_out ),
       .io_VwirePorts_2_20_8_in( ArrayRowModule_2_io_V_wire_out_328 ),
       .io_VwirePorts_2_20_8_en( T1064 ),
       .io_VwirePorts_2_20_8_out( VwireModule_io_VwirePorts_2_20_8_out ),
       .io_VwirePorts_2_20_7_in( ArrayRowModule_2_io_V_wire_out_327 ),
       .io_VwirePorts_2_20_7_en( T1063 ),
       .io_VwirePorts_2_20_7_out( VwireModule_io_VwirePorts_2_20_7_out ),
       .io_VwirePorts_2_20_6_in( ArrayRowModule_2_io_V_wire_out_326 ),
       .io_VwirePorts_2_20_6_en( T1062 ),
       .io_VwirePorts_2_20_6_out( VwireModule_io_VwirePorts_2_20_6_out ),
       .io_VwirePorts_2_20_5_in( ArrayRowModule_2_io_V_wire_out_325 ),
       .io_VwirePorts_2_20_5_en( T1061 ),
       .io_VwirePorts_2_20_5_out( VwireModule_io_VwirePorts_2_20_5_out ),
       .io_VwirePorts_2_20_4_in( ArrayRowModule_2_io_V_wire_out_324 ),
       .io_VwirePorts_2_20_4_en( T1060 ),
       .io_VwirePorts_2_20_4_out( VwireModule_io_VwirePorts_2_20_4_out ),
       .io_VwirePorts_2_20_3_in( ArrayRowModule_2_io_V_wire_out_323 ),
       .io_VwirePorts_2_20_3_en( T1059 ),
       .io_VwirePorts_2_20_3_out( VwireModule_io_VwirePorts_2_20_3_out ),
       .io_VwirePorts_2_20_2_in( ArrayRowModule_2_io_V_wire_out_322 ),
       .io_VwirePorts_2_20_2_en( T1058 ),
       .io_VwirePorts_2_20_2_out( VwireModule_io_VwirePorts_2_20_2_out ),
       .io_VwirePorts_2_20_1_in( ArrayRowModule_2_io_V_wire_out_321 ),
       .io_VwirePorts_2_20_1_en( T1057 ),
       .io_VwirePorts_2_20_1_out( VwireModule_io_VwirePorts_2_20_1_out ),
       .io_VwirePorts_2_20_0_in( ArrayRowModule_2_io_V_wire_out_320 ),
       .io_VwirePorts_2_20_0_en( T1056 ),
       .io_VwirePorts_2_20_0_out( VwireModule_io_VwirePorts_2_20_0_out ),
       .io_VwirePorts_2_19_15_in( ArrayRowModule_2_io_V_wire_out_319 ),
       .io_VwirePorts_2_19_15_en( T1055 ),
       .io_VwirePorts_2_19_15_out( VwireModule_io_VwirePorts_2_19_15_out ),
       .io_VwirePorts_2_19_14_in( ArrayRowModule_2_io_V_wire_out_318 ),
       .io_VwirePorts_2_19_14_en( T1054 ),
       .io_VwirePorts_2_19_14_out( VwireModule_io_VwirePorts_2_19_14_out ),
       .io_VwirePorts_2_19_13_in( ArrayRowModule_2_io_V_wire_out_317 ),
       .io_VwirePorts_2_19_13_en( T1053 ),
       .io_VwirePorts_2_19_13_out( VwireModule_io_VwirePorts_2_19_13_out ),
       .io_VwirePorts_2_19_12_in( ArrayRowModule_2_io_V_wire_out_316 ),
       .io_VwirePorts_2_19_12_en( T1052 ),
       .io_VwirePorts_2_19_12_out( VwireModule_io_VwirePorts_2_19_12_out ),
       .io_VwirePorts_2_19_11_in( ArrayRowModule_2_io_V_wire_out_315 ),
       .io_VwirePorts_2_19_11_en( T1051 ),
       .io_VwirePorts_2_19_11_out( VwireModule_io_VwirePorts_2_19_11_out ),
       .io_VwirePorts_2_19_10_in( ArrayRowModule_2_io_V_wire_out_314 ),
       .io_VwirePorts_2_19_10_en( T1050 ),
       .io_VwirePorts_2_19_10_out( VwireModule_io_VwirePorts_2_19_10_out ),
       .io_VwirePorts_2_19_9_in( ArrayRowModule_2_io_V_wire_out_313 ),
       .io_VwirePorts_2_19_9_en( T1049 ),
       .io_VwirePorts_2_19_9_out( VwireModule_io_VwirePorts_2_19_9_out ),
       .io_VwirePorts_2_19_8_in( ArrayRowModule_2_io_V_wire_out_312 ),
       .io_VwirePorts_2_19_8_en( T1048 ),
       .io_VwirePorts_2_19_8_out( VwireModule_io_VwirePorts_2_19_8_out ),
       .io_VwirePorts_2_19_7_in( ArrayRowModule_2_io_V_wire_out_311 ),
       .io_VwirePorts_2_19_7_en( T1047 ),
       .io_VwirePorts_2_19_7_out( VwireModule_io_VwirePorts_2_19_7_out ),
       .io_VwirePorts_2_19_6_in( ArrayRowModule_2_io_V_wire_out_310 ),
       .io_VwirePorts_2_19_6_en( T1046 ),
       .io_VwirePorts_2_19_6_out( VwireModule_io_VwirePorts_2_19_6_out ),
       .io_VwirePorts_2_19_5_in( ArrayRowModule_2_io_V_wire_out_309 ),
       .io_VwirePorts_2_19_5_en( T1045 ),
       .io_VwirePorts_2_19_5_out( VwireModule_io_VwirePorts_2_19_5_out ),
       .io_VwirePorts_2_19_4_in( ArrayRowModule_2_io_V_wire_out_308 ),
       .io_VwirePorts_2_19_4_en( T1044 ),
       .io_VwirePorts_2_19_4_out( VwireModule_io_VwirePorts_2_19_4_out ),
       .io_VwirePorts_2_19_3_in( ArrayRowModule_2_io_V_wire_out_307 ),
       .io_VwirePorts_2_19_3_en( T1043 ),
       .io_VwirePorts_2_19_3_out( VwireModule_io_VwirePorts_2_19_3_out ),
       .io_VwirePorts_2_19_2_in( ArrayRowModule_2_io_V_wire_out_306 ),
       .io_VwirePorts_2_19_2_en( T1042 ),
       .io_VwirePorts_2_19_2_out( VwireModule_io_VwirePorts_2_19_2_out ),
       .io_VwirePorts_2_19_1_in( ArrayRowModule_2_io_V_wire_out_305 ),
       .io_VwirePorts_2_19_1_en( T1041 ),
       .io_VwirePorts_2_19_1_out( VwireModule_io_VwirePorts_2_19_1_out ),
       .io_VwirePorts_2_19_0_in( ArrayRowModule_2_io_V_wire_out_304 ),
       .io_VwirePorts_2_19_0_en( T1040 ),
       .io_VwirePorts_2_19_0_out( VwireModule_io_VwirePorts_2_19_0_out ),
       .io_VwirePorts_2_18_15_in( ArrayRowModule_2_io_V_wire_out_303 ),
       .io_VwirePorts_2_18_15_en( T1039 ),
       .io_VwirePorts_2_18_15_out( VwireModule_io_VwirePorts_2_18_15_out ),
       .io_VwirePorts_2_18_14_in( ArrayRowModule_2_io_V_wire_out_302 ),
       .io_VwirePorts_2_18_14_en( T1038 ),
       .io_VwirePorts_2_18_14_out( VwireModule_io_VwirePorts_2_18_14_out ),
       .io_VwirePorts_2_18_13_in( ArrayRowModule_2_io_V_wire_out_301 ),
       .io_VwirePorts_2_18_13_en( T1037 ),
       .io_VwirePorts_2_18_13_out( VwireModule_io_VwirePorts_2_18_13_out ),
       .io_VwirePorts_2_18_12_in( ArrayRowModule_2_io_V_wire_out_300 ),
       .io_VwirePorts_2_18_12_en( T1036 ),
       .io_VwirePorts_2_18_12_out( VwireModule_io_VwirePorts_2_18_12_out ),
       .io_VwirePorts_2_18_11_in( ArrayRowModule_2_io_V_wire_out_299 ),
       .io_VwirePorts_2_18_11_en( T1035 ),
       .io_VwirePorts_2_18_11_out( VwireModule_io_VwirePorts_2_18_11_out ),
       .io_VwirePorts_2_18_10_in( ArrayRowModule_2_io_V_wire_out_298 ),
       .io_VwirePorts_2_18_10_en( T1034 ),
       .io_VwirePorts_2_18_10_out( VwireModule_io_VwirePorts_2_18_10_out ),
       .io_VwirePorts_2_18_9_in( ArrayRowModule_2_io_V_wire_out_297 ),
       .io_VwirePorts_2_18_9_en( T1033 ),
       .io_VwirePorts_2_18_9_out( VwireModule_io_VwirePorts_2_18_9_out ),
       .io_VwirePorts_2_18_8_in( ArrayRowModule_2_io_V_wire_out_296 ),
       .io_VwirePorts_2_18_8_en( T1032 ),
       .io_VwirePorts_2_18_8_out( VwireModule_io_VwirePorts_2_18_8_out ),
       .io_VwirePorts_2_18_7_in( ArrayRowModule_2_io_V_wire_out_295 ),
       .io_VwirePorts_2_18_7_en( T1031 ),
       .io_VwirePorts_2_18_7_out( VwireModule_io_VwirePorts_2_18_7_out ),
       .io_VwirePorts_2_18_6_in( ArrayRowModule_2_io_V_wire_out_294 ),
       .io_VwirePorts_2_18_6_en( T1030 ),
       .io_VwirePorts_2_18_6_out( VwireModule_io_VwirePorts_2_18_6_out ),
       .io_VwirePorts_2_18_5_in( ArrayRowModule_2_io_V_wire_out_293 ),
       .io_VwirePorts_2_18_5_en( T1029 ),
       .io_VwirePorts_2_18_5_out( VwireModule_io_VwirePorts_2_18_5_out ),
       .io_VwirePorts_2_18_4_in( ArrayRowModule_2_io_V_wire_out_292 ),
       .io_VwirePorts_2_18_4_en( T1028 ),
       .io_VwirePorts_2_18_4_out( VwireModule_io_VwirePorts_2_18_4_out ),
       .io_VwirePorts_2_18_3_in( ArrayRowModule_2_io_V_wire_out_291 ),
       .io_VwirePorts_2_18_3_en( T1027 ),
       .io_VwirePorts_2_18_3_out( VwireModule_io_VwirePorts_2_18_3_out ),
       .io_VwirePorts_2_18_2_in( ArrayRowModule_2_io_V_wire_out_290 ),
       .io_VwirePorts_2_18_2_en( T1026 ),
       .io_VwirePorts_2_18_2_out( VwireModule_io_VwirePorts_2_18_2_out ),
       .io_VwirePorts_2_18_1_in( ArrayRowModule_2_io_V_wire_out_289 ),
       .io_VwirePorts_2_18_1_en( T1025 ),
       .io_VwirePorts_2_18_1_out( VwireModule_io_VwirePorts_2_18_1_out ),
       .io_VwirePorts_2_18_0_in( ArrayRowModule_2_io_V_wire_out_288 ),
       .io_VwirePorts_2_18_0_en( T1024 ),
       .io_VwirePorts_2_18_0_out( VwireModule_io_VwirePorts_2_18_0_out ),
       .io_VwirePorts_2_17_15_in( ArrayRowModule_2_io_V_wire_out_287 ),
       .io_VwirePorts_2_17_15_en( T1023 ),
       .io_VwirePorts_2_17_15_out( VwireModule_io_VwirePorts_2_17_15_out ),
       .io_VwirePorts_2_17_14_in( ArrayRowModule_2_io_V_wire_out_286 ),
       .io_VwirePorts_2_17_14_en( T1022 ),
       .io_VwirePorts_2_17_14_out( VwireModule_io_VwirePorts_2_17_14_out ),
       .io_VwirePorts_2_17_13_in( ArrayRowModule_2_io_V_wire_out_285 ),
       .io_VwirePorts_2_17_13_en( T1021 ),
       .io_VwirePorts_2_17_13_out( VwireModule_io_VwirePorts_2_17_13_out ),
       .io_VwirePorts_2_17_12_in( ArrayRowModule_2_io_V_wire_out_284 ),
       .io_VwirePorts_2_17_12_en( T1020 ),
       .io_VwirePorts_2_17_12_out( VwireModule_io_VwirePorts_2_17_12_out ),
       .io_VwirePorts_2_17_11_in( ArrayRowModule_2_io_V_wire_out_283 ),
       .io_VwirePorts_2_17_11_en( T1019 ),
       .io_VwirePorts_2_17_11_out( VwireModule_io_VwirePorts_2_17_11_out ),
       .io_VwirePorts_2_17_10_in( ArrayRowModule_2_io_V_wire_out_282 ),
       .io_VwirePorts_2_17_10_en( T1018 ),
       .io_VwirePorts_2_17_10_out( VwireModule_io_VwirePorts_2_17_10_out ),
       .io_VwirePorts_2_17_9_in( ArrayRowModule_2_io_V_wire_out_281 ),
       .io_VwirePorts_2_17_9_en( T1017 ),
       .io_VwirePorts_2_17_9_out( VwireModule_io_VwirePorts_2_17_9_out ),
       .io_VwirePorts_2_17_8_in( ArrayRowModule_2_io_V_wire_out_280 ),
       .io_VwirePorts_2_17_8_en( T1016 ),
       .io_VwirePorts_2_17_8_out( VwireModule_io_VwirePorts_2_17_8_out ),
       .io_VwirePorts_2_17_7_in( ArrayRowModule_2_io_V_wire_out_279 ),
       .io_VwirePorts_2_17_7_en( T1015 ),
       .io_VwirePorts_2_17_7_out( VwireModule_io_VwirePorts_2_17_7_out ),
       .io_VwirePorts_2_17_6_in( ArrayRowModule_2_io_V_wire_out_278 ),
       .io_VwirePorts_2_17_6_en( T1014 ),
       .io_VwirePorts_2_17_6_out( VwireModule_io_VwirePorts_2_17_6_out ),
       .io_VwirePorts_2_17_5_in( ArrayRowModule_2_io_V_wire_out_277 ),
       .io_VwirePorts_2_17_5_en( T1013 ),
       .io_VwirePorts_2_17_5_out( VwireModule_io_VwirePorts_2_17_5_out ),
       .io_VwirePorts_2_17_4_in( ArrayRowModule_2_io_V_wire_out_276 ),
       .io_VwirePorts_2_17_4_en( T1012 ),
       .io_VwirePorts_2_17_4_out( VwireModule_io_VwirePorts_2_17_4_out ),
       .io_VwirePorts_2_17_3_in( ArrayRowModule_2_io_V_wire_out_275 ),
       .io_VwirePorts_2_17_3_en( T1011 ),
       .io_VwirePorts_2_17_3_out( VwireModule_io_VwirePorts_2_17_3_out ),
       .io_VwirePorts_2_17_2_in( ArrayRowModule_2_io_V_wire_out_274 ),
       .io_VwirePorts_2_17_2_en( T1010 ),
       .io_VwirePorts_2_17_2_out( VwireModule_io_VwirePorts_2_17_2_out ),
       .io_VwirePorts_2_17_1_in( ArrayRowModule_2_io_V_wire_out_273 ),
       .io_VwirePorts_2_17_1_en( T1009 ),
       .io_VwirePorts_2_17_1_out( VwireModule_io_VwirePorts_2_17_1_out ),
       .io_VwirePorts_2_17_0_in( ArrayRowModule_2_io_V_wire_out_272 ),
       .io_VwirePorts_2_17_0_en( T1008 ),
       .io_VwirePorts_2_17_0_out( VwireModule_io_VwirePorts_2_17_0_out ),
       .io_VwirePorts_2_16_15_in( ArrayRowModule_2_io_V_wire_out_271 ),
       .io_VwirePorts_2_16_15_en( T1007 ),
       .io_VwirePorts_2_16_15_out( VwireModule_io_VwirePorts_2_16_15_out ),
       .io_VwirePorts_2_16_14_in( ArrayRowModule_2_io_V_wire_out_270 ),
       .io_VwirePorts_2_16_14_en( T1006 ),
       .io_VwirePorts_2_16_14_out( VwireModule_io_VwirePorts_2_16_14_out ),
       .io_VwirePorts_2_16_13_in( ArrayRowModule_2_io_V_wire_out_269 ),
       .io_VwirePorts_2_16_13_en( T1005 ),
       .io_VwirePorts_2_16_13_out( VwireModule_io_VwirePorts_2_16_13_out ),
       .io_VwirePorts_2_16_12_in( ArrayRowModule_2_io_V_wire_out_268 ),
       .io_VwirePorts_2_16_12_en( T1004 ),
       .io_VwirePorts_2_16_12_out( VwireModule_io_VwirePorts_2_16_12_out ),
       .io_VwirePorts_2_16_11_in( ArrayRowModule_2_io_V_wire_out_267 ),
       .io_VwirePorts_2_16_11_en( T1003 ),
       .io_VwirePorts_2_16_11_out( VwireModule_io_VwirePorts_2_16_11_out ),
       .io_VwirePorts_2_16_10_in( ArrayRowModule_2_io_V_wire_out_266 ),
       .io_VwirePorts_2_16_10_en( T1002 ),
       .io_VwirePorts_2_16_10_out( VwireModule_io_VwirePorts_2_16_10_out ),
       .io_VwirePorts_2_16_9_in( ArrayRowModule_2_io_V_wire_out_265 ),
       .io_VwirePorts_2_16_9_en( T1001 ),
       .io_VwirePorts_2_16_9_out( VwireModule_io_VwirePorts_2_16_9_out ),
       .io_VwirePorts_2_16_8_in( ArrayRowModule_2_io_V_wire_out_264 ),
       .io_VwirePorts_2_16_8_en( T1000 ),
       .io_VwirePorts_2_16_8_out( VwireModule_io_VwirePorts_2_16_8_out ),
       .io_VwirePorts_2_16_7_in( ArrayRowModule_2_io_V_wire_out_263 ),
       .io_VwirePorts_2_16_7_en( T999 ),
       .io_VwirePorts_2_16_7_out( VwireModule_io_VwirePorts_2_16_7_out ),
       .io_VwirePorts_2_16_6_in( ArrayRowModule_2_io_V_wire_out_262 ),
       .io_VwirePorts_2_16_6_en( T998 ),
       .io_VwirePorts_2_16_6_out( VwireModule_io_VwirePorts_2_16_6_out ),
       .io_VwirePorts_2_16_5_in( ArrayRowModule_2_io_V_wire_out_261 ),
       .io_VwirePorts_2_16_5_en( T997 ),
       .io_VwirePorts_2_16_5_out( VwireModule_io_VwirePorts_2_16_5_out ),
       .io_VwirePorts_2_16_4_in( ArrayRowModule_2_io_V_wire_out_260 ),
       .io_VwirePorts_2_16_4_en( T996 ),
       .io_VwirePorts_2_16_4_out( VwireModule_io_VwirePorts_2_16_4_out ),
       .io_VwirePorts_2_16_3_in( ArrayRowModule_2_io_V_wire_out_259 ),
       .io_VwirePorts_2_16_3_en( T995 ),
       .io_VwirePorts_2_16_3_out( VwireModule_io_VwirePorts_2_16_3_out ),
       .io_VwirePorts_2_16_2_in( ArrayRowModule_2_io_V_wire_out_258 ),
       .io_VwirePorts_2_16_2_en( T994 ),
       .io_VwirePorts_2_16_2_out( VwireModule_io_VwirePorts_2_16_2_out ),
       .io_VwirePorts_2_16_1_in( ArrayRowModule_2_io_V_wire_out_257 ),
       .io_VwirePorts_2_16_1_en( T993 ),
       .io_VwirePorts_2_16_1_out( VwireModule_io_VwirePorts_2_16_1_out ),
       .io_VwirePorts_2_16_0_in( ArrayRowModule_2_io_V_wire_out_256 ),
       .io_VwirePorts_2_16_0_en( T992 ),
       .io_VwirePorts_2_16_0_out( VwireModule_io_VwirePorts_2_16_0_out ),
       .io_VwirePorts_2_15_15_in( ArrayRowModule_2_io_V_wire_out_255 ),
       .io_VwirePorts_2_15_15_en( T991 ),
       .io_VwirePorts_2_15_15_out( VwireModule_io_VwirePorts_2_15_15_out ),
       .io_VwirePorts_2_15_14_in( ArrayRowModule_2_io_V_wire_out_254 ),
       .io_VwirePorts_2_15_14_en( T990 ),
       .io_VwirePorts_2_15_14_out( VwireModule_io_VwirePorts_2_15_14_out ),
       .io_VwirePorts_2_15_13_in( ArrayRowModule_2_io_V_wire_out_253 ),
       .io_VwirePorts_2_15_13_en( T989 ),
       .io_VwirePorts_2_15_13_out( VwireModule_io_VwirePorts_2_15_13_out ),
       .io_VwirePorts_2_15_12_in( ArrayRowModule_2_io_V_wire_out_252 ),
       .io_VwirePorts_2_15_12_en( T988 ),
       .io_VwirePorts_2_15_12_out( VwireModule_io_VwirePorts_2_15_12_out ),
       .io_VwirePorts_2_15_11_in( ArrayRowModule_2_io_V_wire_out_251 ),
       .io_VwirePorts_2_15_11_en( T987 ),
       .io_VwirePorts_2_15_11_out( VwireModule_io_VwirePorts_2_15_11_out ),
       .io_VwirePorts_2_15_10_in( ArrayRowModule_2_io_V_wire_out_250 ),
       .io_VwirePorts_2_15_10_en( T986 ),
       .io_VwirePorts_2_15_10_out( VwireModule_io_VwirePorts_2_15_10_out ),
       .io_VwirePorts_2_15_9_in( ArrayRowModule_2_io_V_wire_out_249 ),
       .io_VwirePorts_2_15_9_en( T985 ),
       .io_VwirePorts_2_15_9_out( VwireModule_io_VwirePorts_2_15_9_out ),
       .io_VwirePorts_2_15_8_in( ArrayRowModule_2_io_V_wire_out_248 ),
       .io_VwirePorts_2_15_8_en( T984 ),
       .io_VwirePorts_2_15_8_out( VwireModule_io_VwirePorts_2_15_8_out ),
       .io_VwirePorts_2_15_7_in( ArrayRowModule_2_io_V_wire_out_247 ),
       .io_VwirePorts_2_15_7_en( T983 ),
       .io_VwirePorts_2_15_7_out( VwireModule_io_VwirePorts_2_15_7_out ),
       .io_VwirePorts_2_15_6_in( ArrayRowModule_2_io_V_wire_out_246 ),
       .io_VwirePorts_2_15_6_en( T982 ),
       .io_VwirePorts_2_15_6_out( VwireModule_io_VwirePorts_2_15_6_out ),
       .io_VwirePorts_2_15_5_in( ArrayRowModule_2_io_V_wire_out_245 ),
       .io_VwirePorts_2_15_5_en( T981 ),
       .io_VwirePorts_2_15_5_out( VwireModule_io_VwirePorts_2_15_5_out ),
       .io_VwirePorts_2_15_4_in( ArrayRowModule_2_io_V_wire_out_244 ),
       .io_VwirePorts_2_15_4_en( T980 ),
       .io_VwirePorts_2_15_4_out( VwireModule_io_VwirePorts_2_15_4_out ),
       .io_VwirePorts_2_15_3_in( ArrayRowModule_2_io_V_wire_out_243 ),
       .io_VwirePorts_2_15_3_en( T979 ),
       .io_VwirePorts_2_15_3_out( VwireModule_io_VwirePorts_2_15_3_out ),
       .io_VwirePorts_2_15_2_in( ArrayRowModule_2_io_V_wire_out_242 ),
       .io_VwirePorts_2_15_2_en( T978 ),
       .io_VwirePorts_2_15_2_out( VwireModule_io_VwirePorts_2_15_2_out ),
       .io_VwirePorts_2_15_1_in( ArrayRowModule_2_io_V_wire_out_241 ),
       .io_VwirePorts_2_15_1_en( T977 ),
       .io_VwirePorts_2_15_1_out( VwireModule_io_VwirePorts_2_15_1_out ),
       .io_VwirePorts_2_15_0_in( ArrayRowModule_2_io_V_wire_out_240 ),
       .io_VwirePorts_2_15_0_en( T976 ),
       .io_VwirePorts_2_15_0_out( VwireModule_io_VwirePorts_2_15_0_out ),
       .io_VwirePorts_2_14_15_in( ArrayRowModule_2_io_V_wire_out_239 ),
       .io_VwirePorts_2_14_15_en( T975 ),
       .io_VwirePorts_2_14_15_out( VwireModule_io_VwirePorts_2_14_15_out ),
       .io_VwirePorts_2_14_14_in( ArrayRowModule_2_io_V_wire_out_238 ),
       .io_VwirePorts_2_14_14_en( T974 ),
       .io_VwirePorts_2_14_14_out( VwireModule_io_VwirePorts_2_14_14_out ),
       .io_VwirePorts_2_14_13_in( ArrayRowModule_2_io_V_wire_out_237 ),
       .io_VwirePorts_2_14_13_en( T973 ),
       .io_VwirePorts_2_14_13_out( VwireModule_io_VwirePorts_2_14_13_out ),
       .io_VwirePorts_2_14_12_in( ArrayRowModule_2_io_V_wire_out_236 ),
       .io_VwirePorts_2_14_12_en( T972 ),
       .io_VwirePorts_2_14_12_out( VwireModule_io_VwirePorts_2_14_12_out ),
       .io_VwirePorts_2_14_11_in( ArrayRowModule_2_io_V_wire_out_235 ),
       .io_VwirePorts_2_14_11_en( T971 ),
       .io_VwirePorts_2_14_11_out( VwireModule_io_VwirePorts_2_14_11_out ),
       .io_VwirePorts_2_14_10_in( ArrayRowModule_2_io_V_wire_out_234 ),
       .io_VwirePorts_2_14_10_en( T970 ),
       .io_VwirePorts_2_14_10_out( VwireModule_io_VwirePorts_2_14_10_out ),
       .io_VwirePorts_2_14_9_in( ArrayRowModule_2_io_V_wire_out_233 ),
       .io_VwirePorts_2_14_9_en( T969 ),
       .io_VwirePorts_2_14_9_out( VwireModule_io_VwirePorts_2_14_9_out ),
       .io_VwirePorts_2_14_8_in( ArrayRowModule_2_io_V_wire_out_232 ),
       .io_VwirePorts_2_14_8_en( T968 ),
       .io_VwirePorts_2_14_8_out( VwireModule_io_VwirePorts_2_14_8_out ),
       .io_VwirePorts_2_14_7_in( ArrayRowModule_2_io_V_wire_out_231 ),
       .io_VwirePorts_2_14_7_en( T967 ),
       .io_VwirePorts_2_14_7_out( VwireModule_io_VwirePorts_2_14_7_out ),
       .io_VwirePorts_2_14_6_in( ArrayRowModule_2_io_V_wire_out_230 ),
       .io_VwirePorts_2_14_6_en( T966 ),
       .io_VwirePorts_2_14_6_out( VwireModule_io_VwirePorts_2_14_6_out ),
       .io_VwirePorts_2_14_5_in( ArrayRowModule_2_io_V_wire_out_229 ),
       .io_VwirePorts_2_14_5_en( T965 ),
       .io_VwirePorts_2_14_5_out( VwireModule_io_VwirePorts_2_14_5_out ),
       .io_VwirePorts_2_14_4_in( ArrayRowModule_2_io_V_wire_out_228 ),
       .io_VwirePorts_2_14_4_en( T964 ),
       .io_VwirePorts_2_14_4_out( VwireModule_io_VwirePorts_2_14_4_out ),
       .io_VwirePorts_2_14_3_in( ArrayRowModule_2_io_V_wire_out_227 ),
       .io_VwirePorts_2_14_3_en( T963 ),
       .io_VwirePorts_2_14_3_out( VwireModule_io_VwirePorts_2_14_3_out ),
       .io_VwirePorts_2_14_2_in( ArrayRowModule_2_io_V_wire_out_226 ),
       .io_VwirePorts_2_14_2_en( T962 ),
       .io_VwirePorts_2_14_2_out( VwireModule_io_VwirePorts_2_14_2_out ),
       .io_VwirePorts_2_14_1_in( ArrayRowModule_2_io_V_wire_out_225 ),
       .io_VwirePorts_2_14_1_en( T961 ),
       .io_VwirePorts_2_14_1_out( VwireModule_io_VwirePorts_2_14_1_out ),
       .io_VwirePorts_2_14_0_in( ArrayRowModule_2_io_V_wire_out_224 ),
       .io_VwirePorts_2_14_0_en( T960 ),
       .io_VwirePorts_2_14_0_out( VwireModule_io_VwirePorts_2_14_0_out ),
       .io_VwirePorts_2_13_15_in( ArrayRowModule_2_io_V_wire_out_223 ),
       .io_VwirePorts_2_13_15_en( T959 ),
       .io_VwirePorts_2_13_15_out( VwireModule_io_VwirePorts_2_13_15_out ),
       .io_VwirePorts_2_13_14_in( ArrayRowModule_2_io_V_wire_out_222 ),
       .io_VwirePorts_2_13_14_en( T958 ),
       .io_VwirePorts_2_13_14_out( VwireModule_io_VwirePorts_2_13_14_out ),
       .io_VwirePorts_2_13_13_in( ArrayRowModule_2_io_V_wire_out_221 ),
       .io_VwirePorts_2_13_13_en( T957 ),
       .io_VwirePorts_2_13_13_out( VwireModule_io_VwirePorts_2_13_13_out ),
       .io_VwirePorts_2_13_12_in( ArrayRowModule_2_io_V_wire_out_220 ),
       .io_VwirePorts_2_13_12_en( T956 ),
       .io_VwirePorts_2_13_12_out( VwireModule_io_VwirePorts_2_13_12_out ),
       .io_VwirePorts_2_13_11_in( ArrayRowModule_2_io_V_wire_out_219 ),
       .io_VwirePorts_2_13_11_en( T955 ),
       .io_VwirePorts_2_13_11_out( VwireModule_io_VwirePorts_2_13_11_out ),
       .io_VwirePorts_2_13_10_in( ArrayRowModule_2_io_V_wire_out_218 ),
       .io_VwirePorts_2_13_10_en( T954 ),
       .io_VwirePorts_2_13_10_out( VwireModule_io_VwirePorts_2_13_10_out ),
       .io_VwirePorts_2_13_9_in( ArrayRowModule_2_io_V_wire_out_217 ),
       .io_VwirePorts_2_13_9_en( T953 ),
       .io_VwirePorts_2_13_9_out( VwireModule_io_VwirePorts_2_13_9_out ),
       .io_VwirePorts_2_13_8_in( ArrayRowModule_2_io_V_wire_out_216 ),
       .io_VwirePorts_2_13_8_en( T952 ),
       .io_VwirePorts_2_13_8_out( VwireModule_io_VwirePorts_2_13_8_out ),
       .io_VwirePorts_2_13_7_in( ArrayRowModule_2_io_V_wire_out_215 ),
       .io_VwirePorts_2_13_7_en( T951 ),
       .io_VwirePorts_2_13_7_out( VwireModule_io_VwirePorts_2_13_7_out ),
       .io_VwirePorts_2_13_6_in( ArrayRowModule_2_io_V_wire_out_214 ),
       .io_VwirePorts_2_13_6_en( T950 ),
       .io_VwirePorts_2_13_6_out( VwireModule_io_VwirePorts_2_13_6_out ),
       .io_VwirePorts_2_13_5_in( ArrayRowModule_2_io_V_wire_out_213 ),
       .io_VwirePorts_2_13_5_en( T949 ),
       .io_VwirePorts_2_13_5_out( VwireModule_io_VwirePorts_2_13_5_out ),
       .io_VwirePorts_2_13_4_in( ArrayRowModule_2_io_V_wire_out_212 ),
       .io_VwirePorts_2_13_4_en( T948 ),
       .io_VwirePorts_2_13_4_out( VwireModule_io_VwirePorts_2_13_4_out ),
       .io_VwirePorts_2_13_3_in( ArrayRowModule_2_io_V_wire_out_211 ),
       .io_VwirePorts_2_13_3_en( T947 ),
       .io_VwirePorts_2_13_3_out( VwireModule_io_VwirePorts_2_13_3_out ),
       .io_VwirePorts_2_13_2_in( ArrayRowModule_2_io_V_wire_out_210 ),
       .io_VwirePorts_2_13_2_en( T946 ),
       .io_VwirePorts_2_13_2_out( VwireModule_io_VwirePorts_2_13_2_out ),
       .io_VwirePorts_2_13_1_in( ArrayRowModule_2_io_V_wire_out_209 ),
       .io_VwirePorts_2_13_1_en( T945 ),
       .io_VwirePorts_2_13_1_out( VwireModule_io_VwirePorts_2_13_1_out ),
       .io_VwirePorts_2_13_0_in( ArrayRowModule_2_io_V_wire_out_208 ),
       .io_VwirePorts_2_13_0_en( T944 ),
       .io_VwirePorts_2_13_0_out( VwireModule_io_VwirePorts_2_13_0_out ),
       .io_VwirePorts_2_12_15_in( ArrayRowModule_2_io_V_wire_out_207 ),
       .io_VwirePorts_2_12_15_en( T943 ),
       .io_VwirePorts_2_12_15_out( VwireModule_io_VwirePorts_2_12_15_out ),
       .io_VwirePorts_2_12_14_in( ArrayRowModule_2_io_V_wire_out_206 ),
       .io_VwirePorts_2_12_14_en( T942 ),
       .io_VwirePorts_2_12_14_out( VwireModule_io_VwirePorts_2_12_14_out ),
       .io_VwirePorts_2_12_13_in( ArrayRowModule_2_io_V_wire_out_205 ),
       .io_VwirePorts_2_12_13_en( T941 ),
       .io_VwirePorts_2_12_13_out( VwireModule_io_VwirePorts_2_12_13_out ),
       .io_VwirePorts_2_12_12_in( ArrayRowModule_2_io_V_wire_out_204 ),
       .io_VwirePorts_2_12_12_en( T940 ),
       .io_VwirePorts_2_12_12_out( VwireModule_io_VwirePorts_2_12_12_out ),
       .io_VwirePorts_2_12_11_in( ArrayRowModule_2_io_V_wire_out_203 ),
       .io_VwirePorts_2_12_11_en( T939 ),
       .io_VwirePorts_2_12_11_out( VwireModule_io_VwirePorts_2_12_11_out ),
       .io_VwirePorts_2_12_10_in( ArrayRowModule_2_io_V_wire_out_202 ),
       .io_VwirePorts_2_12_10_en( T938 ),
       .io_VwirePorts_2_12_10_out( VwireModule_io_VwirePorts_2_12_10_out ),
       .io_VwirePorts_2_12_9_in( ArrayRowModule_2_io_V_wire_out_201 ),
       .io_VwirePorts_2_12_9_en( T937 ),
       .io_VwirePorts_2_12_9_out( VwireModule_io_VwirePorts_2_12_9_out ),
       .io_VwirePorts_2_12_8_in( ArrayRowModule_2_io_V_wire_out_200 ),
       .io_VwirePorts_2_12_8_en( T936 ),
       .io_VwirePorts_2_12_8_out( VwireModule_io_VwirePorts_2_12_8_out ),
       .io_VwirePorts_2_12_7_in( ArrayRowModule_2_io_V_wire_out_199 ),
       .io_VwirePorts_2_12_7_en( T935 ),
       .io_VwirePorts_2_12_7_out( VwireModule_io_VwirePorts_2_12_7_out ),
       .io_VwirePorts_2_12_6_in( ArrayRowModule_2_io_V_wire_out_198 ),
       .io_VwirePorts_2_12_6_en( T934 ),
       .io_VwirePorts_2_12_6_out( VwireModule_io_VwirePorts_2_12_6_out ),
       .io_VwirePorts_2_12_5_in( ArrayRowModule_2_io_V_wire_out_197 ),
       .io_VwirePorts_2_12_5_en( T933 ),
       .io_VwirePorts_2_12_5_out( VwireModule_io_VwirePorts_2_12_5_out ),
       .io_VwirePorts_2_12_4_in( ArrayRowModule_2_io_V_wire_out_196 ),
       .io_VwirePorts_2_12_4_en( T932 ),
       .io_VwirePorts_2_12_4_out( VwireModule_io_VwirePorts_2_12_4_out ),
       .io_VwirePorts_2_12_3_in( ArrayRowModule_2_io_V_wire_out_195 ),
       .io_VwirePorts_2_12_3_en( T931 ),
       .io_VwirePorts_2_12_3_out( VwireModule_io_VwirePorts_2_12_3_out ),
       .io_VwirePorts_2_12_2_in( ArrayRowModule_2_io_V_wire_out_194 ),
       .io_VwirePorts_2_12_2_en( T930 ),
       .io_VwirePorts_2_12_2_out( VwireModule_io_VwirePorts_2_12_2_out ),
       .io_VwirePorts_2_12_1_in( ArrayRowModule_2_io_V_wire_out_193 ),
       .io_VwirePorts_2_12_1_en( T929 ),
       .io_VwirePorts_2_12_1_out( VwireModule_io_VwirePorts_2_12_1_out ),
       .io_VwirePorts_2_12_0_in( ArrayRowModule_2_io_V_wire_out_192 ),
       .io_VwirePorts_2_12_0_en( T928 ),
       .io_VwirePorts_2_12_0_out( VwireModule_io_VwirePorts_2_12_0_out ),
       .io_VwirePorts_2_11_15_in( ArrayRowModule_2_io_V_wire_out_191 ),
       .io_VwirePorts_2_11_15_en( T927 ),
       .io_VwirePorts_2_11_15_out( VwireModule_io_VwirePorts_2_11_15_out ),
       .io_VwirePorts_2_11_14_in( ArrayRowModule_2_io_V_wire_out_190 ),
       .io_VwirePorts_2_11_14_en( T926 ),
       .io_VwirePorts_2_11_14_out( VwireModule_io_VwirePorts_2_11_14_out ),
       .io_VwirePorts_2_11_13_in( ArrayRowModule_2_io_V_wire_out_189 ),
       .io_VwirePorts_2_11_13_en( T925 ),
       .io_VwirePorts_2_11_13_out( VwireModule_io_VwirePorts_2_11_13_out ),
       .io_VwirePorts_2_11_12_in( ArrayRowModule_2_io_V_wire_out_188 ),
       .io_VwirePorts_2_11_12_en( T924 ),
       .io_VwirePorts_2_11_12_out( VwireModule_io_VwirePorts_2_11_12_out ),
       .io_VwirePorts_2_11_11_in( ArrayRowModule_2_io_V_wire_out_187 ),
       .io_VwirePorts_2_11_11_en( T923 ),
       .io_VwirePorts_2_11_11_out( VwireModule_io_VwirePorts_2_11_11_out ),
       .io_VwirePorts_2_11_10_in( ArrayRowModule_2_io_V_wire_out_186 ),
       .io_VwirePorts_2_11_10_en( T922 ),
       .io_VwirePorts_2_11_10_out( VwireModule_io_VwirePorts_2_11_10_out ),
       .io_VwirePorts_2_11_9_in( ArrayRowModule_2_io_V_wire_out_185 ),
       .io_VwirePorts_2_11_9_en( T921 ),
       .io_VwirePorts_2_11_9_out( VwireModule_io_VwirePorts_2_11_9_out ),
       .io_VwirePorts_2_11_8_in( ArrayRowModule_2_io_V_wire_out_184 ),
       .io_VwirePorts_2_11_8_en( T920 ),
       .io_VwirePorts_2_11_8_out( VwireModule_io_VwirePorts_2_11_8_out ),
       .io_VwirePorts_2_11_7_in( ArrayRowModule_2_io_V_wire_out_183 ),
       .io_VwirePorts_2_11_7_en( T919 ),
       .io_VwirePorts_2_11_7_out( VwireModule_io_VwirePorts_2_11_7_out ),
       .io_VwirePorts_2_11_6_in( ArrayRowModule_2_io_V_wire_out_182 ),
       .io_VwirePorts_2_11_6_en( T918 ),
       .io_VwirePorts_2_11_6_out( VwireModule_io_VwirePorts_2_11_6_out ),
       .io_VwirePorts_2_11_5_in( ArrayRowModule_2_io_V_wire_out_181 ),
       .io_VwirePorts_2_11_5_en( T917 ),
       .io_VwirePorts_2_11_5_out( VwireModule_io_VwirePorts_2_11_5_out ),
       .io_VwirePorts_2_11_4_in( ArrayRowModule_2_io_V_wire_out_180 ),
       .io_VwirePorts_2_11_4_en( T916 ),
       .io_VwirePorts_2_11_4_out( VwireModule_io_VwirePorts_2_11_4_out ),
       .io_VwirePorts_2_11_3_in( ArrayRowModule_2_io_V_wire_out_179 ),
       .io_VwirePorts_2_11_3_en( T915 ),
       .io_VwirePorts_2_11_3_out( VwireModule_io_VwirePorts_2_11_3_out ),
       .io_VwirePorts_2_11_2_in( ArrayRowModule_2_io_V_wire_out_178 ),
       .io_VwirePorts_2_11_2_en( T914 ),
       .io_VwirePorts_2_11_2_out( VwireModule_io_VwirePorts_2_11_2_out ),
       .io_VwirePorts_2_11_1_in( ArrayRowModule_2_io_V_wire_out_177 ),
       .io_VwirePorts_2_11_1_en( T913 ),
       .io_VwirePorts_2_11_1_out( VwireModule_io_VwirePorts_2_11_1_out ),
       .io_VwirePorts_2_11_0_in( ArrayRowModule_2_io_V_wire_out_176 ),
       .io_VwirePorts_2_11_0_en( T912 ),
       .io_VwirePorts_2_11_0_out( VwireModule_io_VwirePorts_2_11_0_out ),
       .io_VwirePorts_2_10_15_in( ArrayRowModule_2_io_V_wire_out_175 ),
       .io_VwirePorts_2_10_15_en( T911 ),
       .io_VwirePorts_2_10_15_out( VwireModule_io_VwirePorts_2_10_15_out ),
       .io_VwirePorts_2_10_14_in( ArrayRowModule_2_io_V_wire_out_174 ),
       .io_VwirePorts_2_10_14_en( T910 ),
       .io_VwirePorts_2_10_14_out( VwireModule_io_VwirePorts_2_10_14_out ),
       .io_VwirePorts_2_10_13_in( ArrayRowModule_2_io_V_wire_out_173 ),
       .io_VwirePorts_2_10_13_en( T909 ),
       .io_VwirePorts_2_10_13_out( VwireModule_io_VwirePorts_2_10_13_out ),
       .io_VwirePorts_2_10_12_in( ArrayRowModule_2_io_V_wire_out_172 ),
       .io_VwirePorts_2_10_12_en( T908 ),
       .io_VwirePorts_2_10_12_out( VwireModule_io_VwirePorts_2_10_12_out ),
       .io_VwirePorts_2_10_11_in( ArrayRowModule_2_io_V_wire_out_171 ),
       .io_VwirePorts_2_10_11_en( T907 ),
       .io_VwirePorts_2_10_11_out( VwireModule_io_VwirePorts_2_10_11_out ),
       .io_VwirePorts_2_10_10_in( ArrayRowModule_2_io_V_wire_out_170 ),
       .io_VwirePorts_2_10_10_en( T906 ),
       .io_VwirePorts_2_10_10_out( VwireModule_io_VwirePorts_2_10_10_out ),
       .io_VwirePorts_2_10_9_in( ArrayRowModule_2_io_V_wire_out_169 ),
       .io_VwirePorts_2_10_9_en( T905 ),
       .io_VwirePorts_2_10_9_out( VwireModule_io_VwirePorts_2_10_9_out ),
       .io_VwirePorts_2_10_8_in( ArrayRowModule_2_io_V_wire_out_168 ),
       .io_VwirePorts_2_10_8_en( T904 ),
       .io_VwirePorts_2_10_8_out( VwireModule_io_VwirePorts_2_10_8_out ),
       .io_VwirePorts_2_10_7_in( ArrayRowModule_2_io_V_wire_out_167 ),
       .io_VwirePorts_2_10_7_en( T903 ),
       .io_VwirePorts_2_10_7_out( VwireModule_io_VwirePorts_2_10_7_out ),
       .io_VwirePorts_2_10_6_in( ArrayRowModule_2_io_V_wire_out_166 ),
       .io_VwirePorts_2_10_6_en( T902 ),
       .io_VwirePorts_2_10_6_out( VwireModule_io_VwirePorts_2_10_6_out ),
       .io_VwirePorts_2_10_5_in( ArrayRowModule_2_io_V_wire_out_165 ),
       .io_VwirePorts_2_10_5_en( T901 ),
       .io_VwirePorts_2_10_5_out( VwireModule_io_VwirePorts_2_10_5_out ),
       .io_VwirePorts_2_10_4_in( ArrayRowModule_2_io_V_wire_out_164 ),
       .io_VwirePorts_2_10_4_en( T900 ),
       .io_VwirePorts_2_10_4_out( VwireModule_io_VwirePorts_2_10_4_out ),
       .io_VwirePorts_2_10_3_in( ArrayRowModule_2_io_V_wire_out_163 ),
       .io_VwirePorts_2_10_3_en( T899 ),
       .io_VwirePorts_2_10_3_out( VwireModule_io_VwirePorts_2_10_3_out ),
       .io_VwirePorts_2_10_2_in( ArrayRowModule_2_io_V_wire_out_162 ),
       .io_VwirePorts_2_10_2_en( T898 ),
       .io_VwirePorts_2_10_2_out( VwireModule_io_VwirePorts_2_10_2_out ),
       .io_VwirePorts_2_10_1_in( ArrayRowModule_2_io_V_wire_out_161 ),
       .io_VwirePorts_2_10_1_en( T897 ),
       .io_VwirePorts_2_10_1_out( VwireModule_io_VwirePorts_2_10_1_out ),
       .io_VwirePorts_2_10_0_in( ArrayRowModule_2_io_V_wire_out_160 ),
       .io_VwirePorts_2_10_0_en( T896 ),
       .io_VwirePorts_2_10_0_out( VwireModule_io_VwirePorts_2_10_0_out ),
       .io_VwirePorts_2_9_15_in( ArrayRowModule_2_io_V_wire_out_159 ),
       .io_VwirePorts_2_9_15_en( T895 ),
       .io_VwirePorts_2_9_15_out( VwireModule_io_VwirePorts_2_9_15_out ),
       .io_VwirePorts_2_9_14_in( ArrayRowModule_2_io_V_wire_out_158 ),
       .io_VwirePorts_2_9_14_en( T894 ),
       .io_VwirePorts_2_9_14_out( VwireModule_io_VwirePorts_2_9_14_out ),
       .io_VwirePorts_2_9_13_in( ArrayRowModule_2_io_V_wire_out_157 ),
       .io_VwirePorts_2_9_13_en( T893 ),
       .io_VwirePorts_2_9_13_out( VwireModule_io_VwirePorts_2_9_13_out ),
       .io_VwirePorts_2_9_12_in( ArrayRowModule_2_io_V_wire_out_156 ),
       .io_VwirePorts_2_9_12_en( T892 ),
       .io_VwirePorts_2_9_12_out( VwireModule_io_VwirePorts_2_9_12_out ),
       .io_VwirePorts_2_9_11_in( ArrayRowModule_2_io_V_wire_out_155 ),
       .io_VwirePorts_2_9_11_en( T891 ),
       .io_VwirePorts_2_9_11_out( VwireModule_io_VwirePorts_2_9_11_out ),
       .io_VwirePorts_2_9_10_in( ArrayRowModule_2_io_V_wire_out_154 ),
       .io_VwirePorts_2_9_10_en( T890 ),
       .io_VwirePorts_2_9_10_out( VwireModule_io_VwirePorts_2_9_10_out ),
       .io_VwirePorts_2_9_9_in( ArrayRowModule_2_io_V_wire_out_153 ),
       .io_VwirePorts_2_9_9_en( T889 ),
       .io_VwirePorts_2_9_9_out( VwireModule_io_VwirePorts_2_9_9_out ),
       .io_VwirePorts_2_9_8_in( ArrayRowModule_2_io_V_wire_out_152 ),
       .io_VwirePorts_2_9_8_en( T888 ),
       .io_VwirePorts_2_9_8_out( VwireModule_io_VwirePorts_2_9_8_out ),
       .io_VwirePorts_2_9_7_in( ArrayRowModule_2_io_V_wire_out_151 ),
       .io_VwirePorts_2_9_7_en( T887 ),
       .io_VwirePorts_2_9_7_out( VwireModule_io_VwirePorts_2_9_7_out ),
       .io_VwirePorts_2_9_6_in( ArrayRowModule_2_io_V_wire_out_150 ),
       .io_VwirePorts_2_9_6_en( T886 ),
       .io_VwirePorts_2_9_6_out( VwireModule_io_VwirePorts_2_9_6_out ),
       .io_VwirePorts_2_9_5_in( ArrayRowModule_2_io_V_wire_out_149 ),
       .io_VwirePorts_2_9_5_en( T885 ),
       .io_VwirePorts_2_9_5_out( VwireModule_io_VwirePorts_2_9_5_out ),
       .io_VwirePorts_2_9_4_in( ArrayRowModule_2_io_V_wire_out_148 ),
       .io_VwirePorts_2_9_4_en( T884 ),
       .io_VwirePorts_2_9_4_out( VwireModule_io_VwirePorts_2_9_4_out ),
       .io_VwirePorts_2_9_3_in( ArrayRowModule_2_io_V_wire_out_147 ),
       .io_VwirePorts_2_9_3_en( T883 ),
       .io_VwirePorts_2_9_3_out( VwireModule_io_VwirePorts_2_9_3_out ),
       .io_VwirePorts_2_9_2_in( ArrayRowModule_2_io_V_wire_out_146 ),
       .io_VwirePorts_2_9_2_en( T882 ),
       .io_VwirePorts_2_9_2_out( VwireModule_io_VwirePorts_2_9_2_out ),
       .io_VwirePorts_2_9_1_in( ArrayRowModule_2_io_V_wire_out_145 ),
       .io_VwirePorts_2_9_1_en( T881 ),
       .io_VwirePorts_2_9_1_out( VwireModule_io_VwirePorts_2_9_1_out ),
       .io_VwirePorts_2_9_0_in( ArrayRowModule_2_io_V_wire_out_144 ),
       .io_VwirePorts_2_9_0_en( T880 ),
       .io_VwirePorts_2_9_0_out( VwireModule_io_VwirePorts_2_9_0_out ),
       .io_VwirePorts_2_8_15_in( ArrayRowModule_2_io_V_wire_out_143 ),
       .io_VwirePorts_2_8_15_en( T879 ),
       .io_VwirePorts_2_8_15_out( VwireModule_io_VwirePorts_2_8_15_out ),
       .io_VwirePorts_2_8_14_in( ArrayRowModule_2_io_V_wire_out_142 ),
       .io_VwirePorts_2_8_14_en( T878 ),
       .io_VwirePorts_2_8_14_out( VwireModule_io_VwirePorts_2_8_14_out ),
       .io_VwirePorts_2_8_13_in( ArrayRowModule_2_io_V_wire_out_141 ),
       .io_VwirePorts_2_8_13_en( T877 ),
       .io_VwirePorts_2_8_13_out( VwireModule_io_VwirePorts_2_8_13_out ),
       .io_VwirePorts_2_8_12_in( ArrayRowModule_2_io_V_wire_out_140 ),
       .io_VwirePorts_2_8_12_en( T876 ),
       .io_VwirePorts_2_8_12_out( VwireModule_io_VwirePorts_2_8_12_out ),
       .io_VwirePorts_2_8_11_in( ArrayRowModule_2_io_V_wire_out_139 ),
       .io_VwirePorts_2_8_11_en( T875 ),
       .io_VwirePorts_2_8_11_out( VwireModule_io_VwirePorts_2_8_11_out ),
       .io_VwirePorts_2_8_10_in( ArrayRowModule_2_io_V_wire_out_138 ),
       .io_VwirePorts_2_8_10_en( T874 ),
       .io_VwirePorts_2_8_10_out( VwireModule_io_VwirePorts_2_8_10_out ),
       .io_VwirePorts_2_8_9_in( ArrayRowModule_2_io_V_wire_out_137 ),
       .io_VwirePorts_2_8_9_en( T873 ),
       .io_VwirePorts_2_8_9_out( VwireModule_io_VwirePorts_2_8_9_out ),
       .io_VwirePorts_2_8_8_in( ArrayRowModule_2_io_V_wire_out_136 ),
       .io_VwirePorts_2_8_8_en( T872 ),
       .io_VwirePorts_2_8_8_out( VwireModule_io_VwirePorts_2_8_8_out ),
       .io_VwirePorts_2_8_7_in( ArrayRowModule_2_io_V_wire_out_135 ),
       .io_VwirePorts_2_8_7_en( T871 ),
       .io_VwirePorts_2_8_7_out( VwireModule_io_VwirePorts_2_8_7_out ),
       .io_VwirePorts_2_8_6_in( ArrayRowModule_2_io_V_wire_out_134 ),
       .io_VwirePorts_2_8_6_en( T870 ),
       .io_VwirePorts_2_8_6_out( VwireModule_io_VwirePorts_2_8_6_out ),
       .io_VwirePorts_2_8_5_in( ArrayRowModule_2_io_V_wire_out_133 ),
       .io_VwirePorts_2_8_5_en( T869 ),
       .io_VwirePorts_2_8_5_out( VwireModule_io_VwirePorts_2_8_5_out ),
       .io_VwirePorts_2_8_4_in( ArrayRowModule_2_io_V_wire_out_132 ),
       .io_VwirePorts_2_8_4_en( T868 ),
       .io_VwirePorts_2_8_4_out( VwireModule_io_VwirePorts_2_8_4_out ),
       .io_VwirePorts_2_8_3_in( ArrayRowModule_2_io_V_wire_out_131 ),
       .io_VwirePorts_2_8_3_en( T867 ),
       .io_VwirePorts_2_8_3_out( VwireModule_io_VwirePorts_2_8_3_out ),
       .io_VwirePorts_2_8_2_in( ArrayRowModule_2_io_V_wire_out_130 ),
       .io_VwirePorts_2_8_2_en( T866 ),
       .io_VwirePorts_2_8_2_out( VwireModule_io_VwirePorts_2_8_2_out ),
       .io_VwirePorts_2_8_1_in( ArrayRowModule_2_io_V_wire_out_129 ),
       .io_VwirePorts_2_8_1_en( T865 ),
       .io_VwirePorts_2_8_1_out( VwireModule_io_VwirePorts_2_8_1_out ),
       .io_VwirePorts_2_8_0_in( ArrayRowModule_2_io_V_wire_out_128 ),
       .io_VwirePorts_2_8_0_en( T864 ),
       .io_VwirePorts_2_8_0_out( VwireModule_io_VwirePorts_2_8_0_out ),
       .io_VwirePorts_2_7_15_in( ArrayRowModule_2_io_V_wire_out_127 ),
       .io_VwirePorts_2_7_15_en( T863 ),
       .io_VwirePorts_2_7_15_out( VwireModule_io_VwirePorts_2_7_15_out ),
       .io_VwirePorts_2_7_14_in( ArrayRowModule_2_io_V_wire_out_126 ),
       .io_VwirePorts_2_7_14_en( T862 ),
       .io_VwirePorts_2_7_14_out( VwireModule_io_VwirePorts_2_7_14_out ),
       .io_VwirePorts_2_7_13_in( ArrayRowModule_2_io_V_wire_out_125 ),
       .io_VwirePorts_2_7_13_en( T861 ),
       .io_VwirePorts_2_7_13_out( VwireModule_io_VwirePorts_2_7_13_out ),
       .io_VwirePorts_2_7_12_in( ArrayRowModule_2_io_V_wire_out_124 ),
       .io_VwirePorts_2_7_12_en( T860 ),
       .io_VwirePorts_2_7_12_out( VwireModule_io_VwirePorts_2_7_12_out ),
       .io_VwirePorts_2_7_11_in( ArrayRowModule_2_io_V_wire_out_123 ),
       .io_VwirePorts_2_7_11_en( T859 ),
       .io_VwirePorts_2_7_11_out( VwireModule_io_VwirePorts_2_7_11_out ),
       .io_VwirePorts_2_7_10_in( ArrayRowModule_2_io_V_wire_out_122 ),
       .io_VwirePorts_2_7_10_en( T858 ),
       .io_VwirePorts_2_7_10_out( VwireModule_io_VwirePorts_2_7_10_out ),
       .io_VwirePorts_2_7_9_in( ArrayRowModule_2_io_V_wire_out_121 ),
       .io_VwirePorts_2_7_9_en( T857 ),
       .io_VwirePorts_2_7_9_out( VwireModule_io_VwirePorts_2_7_9_out ),
       .io_VwirePorts_2_7_8_in( ArrayRowModule_2_io_V_wire_out_120 ),
       .io_VwirePorts_2_7_8_en( T856 ),
       .io_VwirePorts_2_7_8_out( VwireModule_io_VwirePorts_2_7_8_out ),
       .io_VwirePorts_2_7_7_in( ArrayRowModule_2_io_V_wire_out_119 ),
       .io_VwirePorts_2_7_7_en( T855 ),
       .io_VwirePorts_2_7_7_out( VwireModule_io_VwirePorts_2_7_7_out ),
       .io_VwirePorts_2_7_6_in( ArrayRowModule_2_io_V_wire_out_118 ),
       .io_VwirePorts_2_7_6_en( T854 ),
       .io_VwirePorts_2_7_6_out( VwireModule_io_VwirePorts_2_7_6_out ),
       .io_VwirePorts_2_7_5_in( ArrayRowModule_2_io_V_wire_out_117 ),
       .io_VwirePorts_2_7_5_en( T853 ),
       .io_VwirePorts_2_7_5_out( VwireModule_io_VwirePorts_2_7_5_out ),
       .io_VwirePorts_2_7_4_in( ArrayRowModule_2_io_V_wire_out_116 ),
       .io_VwirePorts_2_7_4_en( T852 ),
       .io_VwirePorts_2_7_4_out( VwireModule_io_VwirePorts_2_7_4_out ),
       .io_VwirePorts_2_7_3_in( ArrayRowModule_2_io_V_wire_out_115 ),
       .io_VwirePorts_2_7_3_en( T851 ),
       .io_VwirePorts_2_7_3_out( VwireModule_io_VwirePorts_2_7_3_out ),
       .io_VwirePorts_2_7_2_in( ArrayRowModule_2_io_V_wire_out_114 ),
       .io_VwirePorts_2_7_2_en( T850 ),
       .io_VwirePorts_2_7_2_out( VwireModule_io_VwirePorts_2_7_2_out ),
       .io_VwirePorts_2_7_1_in( ArrayRowModule_2_io_V_wire_out_113 ),
       .io_VwirePorts_2_7_1_en( T849 ),
       .io_VwirePorts_2_7_1_out( VwireModule_io_VwirePorts_2_7_1_out ),
       .io_VwirePorts_2_7_0_in( ArrayRowModule_2_io_V_wire_out_112 ),
       .io_VwirePorts_2_7_0_en( T848 ),
       .io_VwirePorts_2_7_0_out( VwireModule_io_VwirePorts_2_7_0_out ),
       .io_VwirePorts_2_6_15_in( ArrayRowModule_2_io_V_wire_out_111 ),
       .io_VwirePorts_2_6_15_en( T847 ),
       .io_VwirePorts_2_6_15_out( VwireModule_io_VwirePorts_2_6_15_out ),
       .io_VwirePorts_2_6_14_in( ArrayRowModule_2_io_V_wire_out_110 ),
       .io_VwirePorts_2_6_14_en( T846 ),
       .io_VwirePorts_2_6_14_out( VwireModule_io_VwirePorts_2_6_14_out ),
       .io_VwirePorts_2_6_13_in( ArrayRowModule_2_io_V_wire_out_109 ),
       .io_VwirePorts_2_6_13_en( T845 ),
       .io_VwirePorts_2_6_13_out( VwireModule_io_VwirePorts_2_6_13_out ),
       .io_VwirePorts_2_6_12_in( ArrayRowModule_2_io_V_wire_out_108 ),
       .io_VwirePorts_2_6_12_en( T844 ),
       .io_VwirePorts_2_6_12_out( VwireModule_io_VwirePorts_2_6_12_out ),
       .io_VwirePorts_2_6_11_in( ArrayRowModule_2_io_V_wire_out_107 ),
       .io_VwirePorts_2_6_11_en( T843 ),
       .io_VwirePorts_2_6_11_out( VwireModule_io_VwirePorts_2_6_11_out ),
       .io_VwirePorts_2_6_10_in( ArrayRowModule_2_io_V_wire_out_106 ),
       .io_VwirePorts_2_6_10_en( T842 ),
       .io_VwirePorts_2_6_10_out( VwireModule_io_VwirePorts_2_6_10_out ),
       .io_VwirePorts_2_6_9_in( ArrayRowModule_2_io_V_wire_out_105 ),
       .io_VwirePorts_2_6_9_en( T841 ),
       .io_VwirePorts_2_6_9_out( VwireModule_io_VwirePorts_2_6_9_out ),
       .io_VwirePorts_2_6_8_in( ArrayRowModule_2_io_V_wire_out_104 ),
       .io_VwirePorts_2_6_8_en( T840 ),
       .io_VwirePorts_2_6_8_out( VwireModule_io_VwirePorts_2_6_8_out ),
       .io_VwirePorts_2_6_7_in( ArrayRowModule_2_io_V_wire_out_103 ),
       .io_VwirePorts_2_6_7_en( T839 ),
       .io_VwirePorts_2_6_7_out( VwireModule_io_VwirePorts_2_6_7_out ),
       .io_VwirePorts_2_6_6_in( ArrayRowModule_2_io_V_wire_out_102 ),
       .io_VwirePorts_2_6_6_en( T838 ),
       .io_VwirePorts_2_6_6_out( VwireModule_io_VwirePorts_2_6_6_out ),
       .io_VwirePorts_2_6_5_in( ArrayRowModule_2_io_V_wire_out_101 ),
       .io_VwirePorts_2_6_5_en( T837 ),
       .io_VwirePorts_2_6_5_out( VwireModule_io_VwirePorts_2_6_5_out ),
       .io_VwirePorts_2_6_4_in( ArrayRowModule_2_io_V_wire_out_100 ),
       .io_VwirePorts_2_6_4_en( T836 ),
       .io_VwirePorts_2_6_4_out( VwireModule_io_VwirePorts_2_6_4_out ),
       .io_VwirePorts_2_6_3_in( ArrayRowModule_2_io_V_wire_out_99 ),
       .io_VwirePorts_2_6_3_en( T835 ),
       .io_VwirePorts_2_6_3_out( VwireModule_io_VwirePorts_2_6_3_out ),
       .io_VwirePorts_2_6_2_in( ArrayRowModule_2_io_V_wire_out_98 ),
       .io_VwirePorts_2_6_2_en( T834 ),
       .io_VwirePorts_2_6_2_out( VwireModule_io_VwirePorts_2_6_2_out ),
       .io_VwirePorts_2_6_1_in( ArrayRowModule_2_io_V_wire_out_97 ),
       .io_VwirePorts_2_6_1_en( T833 ),
       .io_VwirePorts_2_6_1_out( VwireModule_io_VwirePorts_2_6_1_out ),
       .io_VwirePorts_2_6_0_in( ArrayRowModule_2_io_V_wire_out_96 ),
       .io_VwirePorts_2_6_0_en( T832 ),
       .io_VwirePorts_2_6_0_out( VwireModule_io_VwirePorts_2_6_0_out ),
       .io_VwirePorts_2_5_15_in( ArrayRowModule_2_io_V_wire_out_95 ),
       .io_VwirePorts_2_5_15_en( T831 ),
       .io_VwirePorts_2_5_15_out( VwireModule_io_VwirePorts_2_5_15_out ),
       .io_VwirePorts_2_5_14_in( ArrayRowModule_2_io_V_wire_out_94 ),
       .io_VwirePorts_2_5_14_en( T830 ),
       .io_VwirePorts_2_5_14_out( VwireModule_io_VwirePorts_2_5_14_out ),
       .io_VwirePorts_2_5_13_in( ArrayRowModule_2_io_V_wire_out_93 ),
       .io_VwirePorts_2_5_13_en( T829 ),
       .io_VwirePorts_2_5_13_out( VwireModule_io_VwirePorts_2_5_13_out ),
       .io_VwirePorts_2_5_12_in( ArrayRowModule_2_io_V_wire_out_92 ),
       .io_VwirePorts_2_5_12_en( T828 ),
       .io_VwirePorts_2_5_12_out( VwireModule_io_VwirePorts_2_5_12_out ),
       .io_VwirePorts_2_5_11_in( ArrayRowModule_2_io_V_wire_out_91 ),
       .io_VwirePorts_2_5_11_en( T827 ),
       .io_VwirePorts_2_5_11_out( VwireModule_io_VwirePorts_2_5_11_out ),
       .io_VwirePorts_2_5_10_in( ArrayRowModule_2_io_V_wire_out_90 ),
       .io_VwirePorts_2_5_10_en( T826 ),
       .io_VwirePorts_2_5_10_out( VwireModule_io_VwirePorts_2_5_10_out ),
       .io_VwirePorts_2_5_9_in( ArrayRowModule_2_io_V_wire_out_89 ),
       .io_VwirePorts_2_5_9_en( T825 ),
       .io_VwirePorts_2_5_9_out( VwireModule_io_VwirePorts_2_5_9_out ),
       .io_VwirePorts_2_5_8_in( ArrayRowModule_2_io_V_wire_out_88 ),
       .io_VwirePorts_2_5_8_en( T824 ),
       .io_VwirePorts_2_5_8_out( VwireModule_io_VwirePorts_2_5_8_out ),
       .io_VwirePorts_2_5_7_in( ArrayRowModule_2_io_V_wire_out_87 ),
       .io_VwirePorts_2_5_7_en( T823 ),
       .io_VwirePorts_2_5_7_out( VwireModule_io_VwirePorts_2_5_7_out ),
       .io_VwirePorts_2_5_6_in( ArrayRowModule_2_io_V_wire_out_86 ),
       .io_VwirePorts_2_5_6_en( T822 ),
       .io_VwirePorts_2_5_6_out( VwireModule_io_VwirePorts_2_5_6_out ),
       .io_VwirePorts_2_5_5_in( ArrayRowModule_2_io_V_wire_out_85 ),
       .io_VwirePorts_2_5_5_en( T821 ),
       .io_VwirePorts_2_5_5_out( VwireModule_io_VwirePorts_2_5_5_out ),
       .io_VwirePorts_2_5_4_in( ArrayRowModule_2_io_V_wire_out_84 ),
       .io_VwirePorts_2_5_4_en( T820 ),
       .io_VwirePorts_2_5_4_out( VwireModule_io_VwirePorts_2_5_4_out ),
       .io_VwirePorts_2_5_3_in( ArrayRowModule_2_io_V_wire_out_83 ),
       .io_VwirePorts_2_5_3_en( T819 ),
       .io_VwirePorts_2_5_3_out( VwireModule_io_VwirePorts_2_5_3_out ),
       .io_VwirePorts_2_5_2_in( ArrayRowModule_2_io_V_wire_out_82 ),
       .io_VwirePorts_2_5_2_en( T818 ),
       .io_VwirePorts_2_5_2_out( VwireModule_io_VwirePorts_2_5_2_out ),
       .io_VwirePorts_2_5_1_in( ArrayRowModule_2_io_V_wire_out_81 ),
       .io_VwirePorts_2_5_1_en( T817 ),
       .io_VwirePorts_2_5_1_out( VwireModule_io_VwirePorts_2_5_1_out ),
       .io_VwirePorts_2_5_0_in( ArrayRowModule_2_io_V_wire_out_80 ),
       .io_VwirePorts_2_5_0_en( T816 ),
       .io_VwirePorts_2_5_0_out( VwireModule_io_VwirePorts_2_5_0_out ),
       .io_VwirePorts_2_4_15_in( ArrayRowModule_2_io_V_wire_out_79 ),
       .io_VwirePorts_2_4_15_en( T815 ),
       .io_VwirePorts_2_4_15_out( VwireModule_io_VwirePorts_2_4_15_out ),
       .io_VwirePorts_2_4_14_in( ArrayRowModule_2_io_V_wire_out_78 ),
       .io_VwirePorts_2_4_14_en( T814 ),
       .io_VwirePorts_2_4_14_out( VwireModule_io_VwirePorts_2_4_14_out ),
       .io_VwirePorts_2_4_13_in( ArrayRowModule_2_io_V_wire_out_77 ),
       .io_VwirePorts_2_4_13_en( T813 ),
       .io_VwirePorts_2_4_13_out( VwireModule_io_VwirePorts_2_4_13_out ),
       .io_VwirePorts_2_4_12_in( ArrayRowModule_2_io_V_wire_out_76 ),
       .io_VwirePorts_2_4_12_en( T812 ),
       .io_VwirePorts_2_4_12_out( VwireModule_io_VwirePorts_2_4_12_out ),
       .io_VwirePorts_2_4_11_in( ArrayRowModule_2_io_V_wire_out_75 ),
       .io_VwirePorts_2_4_11_en( T811 ),
       .io_VwirePorts_2_4_11_out( VwireModule_io_VwirePorts_2_4_11_out ),
       .io_VwirePorts_2_4_10_in( ArrayRowModule_2_io_V_wire_out_74 ),
       .io_VwirePorts_2_4_10_en( T810 ),
       .io_VwirePorts_2_4_10_out( VwireModule_io_VwirePorts_2_4_10_out ),
       .io_VwirePorts_2_4_9_in( ArrayRowModule_2_io_V_wire_out_73 ),
       .io_VwirePorts_2_4_9_en( T809 ),
       .io_VwirePorts_2_4_9_out( VwireModule_io_VwirePorts_2_4_9_out ),
       .io_VwirePorts_2_4_8_in( ArrayRowModule_2_io_V_wire_out_72 ),
       .io_VwirePorts_2_4_8_en( T808 ),
       .io_VwirePorts_2_4_8_out( VwireModule_io_VwirePorts_2_4_8_out ),
       .io_VwirePorts_2_4_7_in( ArrayRowModule_2_io_V_wire_out_71 ),
       .io_VwirePorts_2_4_7_en( T807 ),
       .io_VwirePorts_2_4_7_out( VwireModule_io_VwirePorts_2_4_7_out ),
       .io_VwirePorts_2_4_6_in( ArrayRowModule_2_io_V_wire_out_70 ),
       .io_VwirePorts_2_4_6_en( T806 ),
       .io_VwirePorts_2_4_6_out( VwireModule_io_VwirePorts_2_4_6_out ),
       .io_VwirePorts_2_4_5_in( ArrayRowModule_2_io_V_wire_out_69 ),
       .io_VwirePorts_2_4_5_en( T805 ),
       .io_VwirePorts_2_4_5_out( VwireModule_io_VwirePorts_2_4_5_out ),
       .io_VwirePorts_2_4_4_in( ArrayRowModule_2_io_V_wire_out_68 ),
       .io_VwirePorts_2_4_4_en( T804 ),
       .io_VwirePorts_2_4_4_out( VwireModule_io_VwirePorts_2_4_4_out ),
       .io_VwirePorts_2_4_3_in( ArrayRowModule_2_io_V_wire_out_67 ),
       .io_VwirePorts_2_4_3_en( T803 ),
       .io_VwirePorts_2_4_3_out( VwireModule_io_VwirePorts_2_4_3_out ),
       .io_VwirePorts_2_4_2_in( ArrayRowModule_2_io_V_wire_out_66 ),
       .io_VwirePorts_2_4_2_en( T802 ),
       .io_VwirePorts_2_4_2_out( VwireModule_io_VwirePorts_2_4_2_out ),
       .io_VwirePorts_2_4_1_in( ArrayRowModule_2_io_V_wire_out_65 ),
       .io_VwirePorts_2_4_1_en( T801 ),
       .io_VwirePorts_2_4_1_out( VwireModule_io_VwirePorts_2_4_1_out ),
       .io_VwirePorts_2_4_0_in( ArrayRowModule_2_io_V_wire_out_64 ),
       .io_VwirePorts_2_4_0_en( T800 ),
       .io_VwirePorts_2_4_0_out( VwireModule_io_VwirePorts_2_4_0_out ),
       .io_VwirePorts_2_3_15_in( ArrayRowModule_2_io_V_wire_out_63 ),
       .io_VwirePorts_2_3_15_en( T799 ),
       .io_VwirePorts_2_3_15_out( VwireModule_io_VwirePorts_2_3_15_out ),
       .io_VwirePorts_2_3_14_in( ArrayRowModule_2_io_V_wire_out_62 ),
       .io_VwirePorts_2_3_14_en( T798 ),
       .io_VwirePorts_2_3_14_out( VwireModule_io_VwirePorts_2_3_14_out ),
       .io_VwirePorts_2_3_13_in( ArrayRowModule_2_io_V_wire_out_61 ),
       .io_VwirePorts_2_3_13_en( T797 ),
       .io_VwirePorts_2_3_13_out( VwireModule_io_VwirePorts_2_3_13_out ),
       .io_VwirePorts_2_3_12_in( ArrayRowModule_2_io_V_wire_out_60 ),
       .io_VwirePorts_2_3_12_en( T796 ),
       .io_VwirePorts_2_3_12_out( VwireModule_io_VwirePorts_2_3_12_out ),
       .io_VwirePorts_2_3_11_in( ArrayRowModule_2_io_V_wire_out_59 ),
       .io_VwirePorts_2_3_11_en( T795 ),
       .io_VwirePorts_2_3_11_out( VwireModule_io_VwirePorts_2_3_11_out ),
       .io_VwirePorts_2_3_10_in( ArrayRowModule_2_io_V_wire_out_58 ),
       .io_VwirePorts_2_3_10_en( T794 ),
       .io_VwirePorts_2_3_10_out( VwireModule_io_VwirePorts_2_3_10_out ),
       .io_VwirePorts_2_3_9_in( ArrayRowModule_2_io_V_wire_out_57 ),
       .io_VwirePorts_2_3_9_en( T793 ),
       .io_VwirePorts_2_3_9_out( VwireModule_io_VwirePorts_2_3_9_out ),
       .io_VwirePorts_2_3_8_in( ArrayRowModule_2_io_V_wire_out_56 ),
       .io_VwirePorts_2_3_8_en( T792 ),
       .io_VwirePorts_2_3_8_out( VwireModule_io_VwirePorts_2_3_8_out ),
       .io_VwirePorts_2_3_7_in( ArrayRowModule_2_io_V_wire_out_55 ),
       .io_VwirePorts_2_3_7_en( T791 ),
       .io_VwirePorts_2_3_7_out( VwireModule_io_VwirePorts_2_3_7_out ),
       .io_VwirePorts_2_3_6_in( ArrayRowModule_2_io_V_wire_out_54 ),
       .io_VwirePorts_2_3_6_en( T790 ),
       .io_VwirePorts_2_3_6_out( VwireModule_io_VwirePorts_2_3_6_out ),
       .io_VwirePorts_2_3_5_in( ArrayRowModule_2_io_V_wire_out_53 ),
       .io_VwirePorts_2_3_5_en( T789 ),
       .io_VwirePorts_2_3_5_out( VwireModule_io_VwirePorts_2_3_5_out ),
       .io_VwirePorts_2_3_4_in( ArrayRowModule_2_io_V_wire_out_52 ),
       .io_VwirePorts_2_3_4_en( T788 ),
       .io_VwirePorts_2_3_4_out( VwireModule_io_VwirePorts_2_3_4_out ),
       .io_VwirePorts_2_3_3_in( ArrayRowModule_2_io_V_wire_out_51 ),
       .io_VwirePorts_2_3_3_en( T787 ),
       .io_VwirePorts_2_3_3_out( VwireModule_io_VwirePorts_2_3_3_out ),
       .io_VwirePorts_2_3_2_in( ArrayRowModule_2_io_V_wire_out_50 ),
       .io_VwirePorts_2_3_2_en( T786 ),
       .io_VwirePorts_2_3_2_out( VwireModule_io_VwirePorts_2_3_2_out ),
       .io_VwirePorts_2_3_1_in( ArrayRowModule_2_io_V_wire_out_49 ),
       .io_VwirePorts_2_3_1_en( T785 ),
       .io_VwirePorts_2_3_1_out( VwireModule_io_VwirePorts_2_3_1_out ),
       .io_VwirePorts_2_3_0_in( ArrayRowModule_2_io_V_wire_out_48 ),
       .io_VwirePorts_2_3_0_en( T784 ),
       .io_VwirePorts_2_3_0_out( VwireModule_io_VwirePorts_2_3_0_out ),
       .io_VwirePorts_2_2_15_in( ArrayRowModule_2_io_V_wire_out_47 ),
       .io_VwirePorts_2_2_15_en( T783 ),
       .io_VwirePorts_2_2_15_out( VwireModule_io_VwirePorts_2_2_15_out ),
       .io_VwirePorts_2_2_14_in( ArrayRowModule_2_io_V_wire_out_46 ),
       .io_VwirePorts_2_2_14_en( T782 ),
       .io_VwirePorts_2_2_14_out( VwireModule_io_VwirePorts_2_2_14_out ),
       .io_VwirePorts_2_2_13_in( ArrayRowModule_2_io_V_wire_out_45 ),
       .io_VwirePorts_2_2_13_en( T781 ),
       .io_VwirePorts_2_2_13_out( VwireModule_io_VwirePorts_2_2_13_out ),
       .io_VwirePorts_2_2_12_in( ArrayRowModule_2_io_V_wire_out_44 ),
       .io_VwirePorts_2_2_12_en( T780 ),
       .io_VwirePorts_2_2_12_out( VwireModule_io_VwirePorts_2_2_12_out ),
       .io_VwirePorts_2_2_11_in( ArrayRowModule_2_io_V_wire_out_43 ),
       .io_VwirePorts_2_2_11_en( T779 ),
       .io_VwirePorts_2_2_11_out( VwireModule_io_VwirePorts_2_2_11_out ),
       .io_VwirePorts_2_2_10_in( ArrayRowModule_2_io_V_wire_out_42 ),
       .io_VwirePorts_2_2_10_en( T778 ),
       .io_VwirePorts_2_2_10_out( VwireModule_io_VwirePorts_2_2_10_out ),
       .io_VwirePorts_2_2_9_in( ArrayRowModule_2_io_V_wire_out_41 ),
       .io_VwirePorts_2_2_9_en( T777 ),
       .io_VwirePorts_2_2_9_out( VwireModule_io_VwirePorts_2_2_9_out ),
       .io_VwirePorts_2_2_8_in( ArrayRowModule_2_io_V_wire_out_40 ),
       .io_VwirePorts_2_2_8_en( T776 ),
       .io_VwirePorts_2_2_8_out( VwireModule_io_VwirePorts_2_2_8_out ),
       .io_VwirePorts_2_2_7_in( ArrayRowModule_2_io_V_wire_out_39 ),
       .io_VwirePorts_2_2_7_en( T775 ),
       .io_VwirePorts_2_2_7_out( VwireModule_io_VwirePorts_2_2_7_out ),
       .io_VwirePorts_2_2_6_in( ArrayRowModule_2_io_V_wire_out_38 ),
       .io_VwirePorts_2_2_6_en( T774 ),
       .io_VwirePorts_2_2_6_out( VwireModule_io_VwirePorts_2_2_6_out ),
       .io_VwirePorts_2_2_5_in( ArrayRowModule_2_io_V_wire_out_37 ),
       .io_VwirePorts_2_2_5_en( T773 ),
       .io_VwirePorts_2_2_5_out( VwireModule_io_VwirePorts_2_2_5_out ),
       .io_VwirePorts_2_2_4_in( ArrayRowModule_2_io_V_wire_out_36 ),
       .io_VwirePorts_2_2_4_en( T772 ),
       .io_VwirePorts_2_2_4_out( VwireModule_io_VwirePorts_2_2_4_out ),
       .io_VwirePorts_2_2_3_in( ArrayRowModule_2_io_V_wire_out_35 ),
       .io_VwirePorts_2_2_3_en( T771 ),
       .io_VwirePorts_2_2_3_out( VwireModule_io_VwirePorts_2_2_3_out ),
       .io_VwirePorts_2_2_2_in( ArrayRowModule_2_io_V_wire_out_34 ),
       .io_VwirePorts_2_2_2_en( T770 ),
       .io_VwirePorts_2_2_2_out( VwireModule_io_VwirePorts_2_2_2_out ),
       .io_VwirePorts_2_2_1_in( ArrayRowModule_2_io_V_wire_out_33 ),
       .io_VwirePorts_2_2_1_en( T769 ),
       .io_VwirePorts_2_2_1_out( VwireModule_io_VwirePorts_2_2_1_out ),
       .io_VwirePorts_2_2_0_in( ArrayRowModule_2_io_V_wire_out_32 ),
       .io_VwirePorts_2_2_0_en( T768 ),
       .io_VwirePorts_2_2_0_out( VwireModule_io_VwirePorts_2_2_0_out ),
       .io_VwirePorts_2_1_15_in( ArrayRowModule_2_io_V_wire_out_31 ),
       .io_VwirePorts_2_1_15_en( T767 ),
       .io_VwirePorts_2_1_15_out( VwireModule_io_VwirePorts_2_1_15_out ),
       .io_VwirePorts_2_1_14_in( ArrayRowModule_2_io_V_wire_out_30 ),
       .io_VwirePorts_2_1_14_en( T766 ),
       .io_VwirePorts_2_1_14_out( VwireModule_io_VwirePorts_2_1_14_out ),
       .io_VwirePorts_2_1_13_in( ArrayRowModule_2_io_V_wire_out_29 ),
       .io_VwirePorts_2_1_13_en( T765 ),
       .io_VwirePorts_2_1_13_out( VwireModule_io_VwirePorts_2_1_13_out ),
       .io_VwirePorts_2_1_12_in( ArrayRowModule_2_io_V_wire_out_28 ),
       .io_VwirePorts_2_1_12_en( T764 ),
       .io_VwirePorts_2_1_12_out( VwireModule_io_VwirePorts_2_1_12_out ),
       .io_VwirePorts_2_1_11_in( ArrayRowModule_2_io_V_wire_out_27 ),
       .io_VwirePorts_2_1_11_en( T763 ),
       .io_VwirePorts_2_1_11_out( VwireModule_io_VwirePorts_2_1_11_out ),
       .io_VwirePorts_2_1_10_in( ArrayRowModule_2_io_V_wire_out_26 ),
       .io_VwirePorts_2_1_10_en( T762 ),
       .io_VwirePorts_2_1_10_out( VwireModule_io_VwirePorts_2_1_10_out ),
       .io_VwirePorts_2_1_9_in( ArrayRowModule_2_io_V_wire_out_25 ),
       .io_VwirePorts_2_1_9_en( T761 ),
       .io_VwirePorts_2_1_9_out( VwireModule_io_VwirePorts_2_1_9_out ),
       .io_VwirePorts_2_1_8_in( ArrayRowModule_2_io_V_wire_out_24 ),
       .io_VwirePorts_2_1_8_en( T760 ),
       .io_VwirePorts_2_1_8_out( VwireModule_io_VwirePorts_2_1_8_out ),
       .io_VwirePorts_2_1_7_in( ArrayRowModule_2_io_V_wire_out_23 ),
       .io_VwirePorts_2_1_7_en( T759 ),
       .io_VwirePorts_2_1_7_out( VwireModule_io_VwirePorts_2_1_7_out ),
       .io_VwirePorts_2_1_6_in( ArrayRowModule_2_io_V_wire_out_22 ),
       .io_VwirePorts_2_1_6_en( T758 ),
       .io_VwirePorts_2_1_6_out( VwireModule_io_VwirePorts_2_1_6_out ),
       .io_VwirePorts_2_1_5_in( ArrayRowModule_2_io_V_wire_out_21 ),
       .io_VwirePorts_2_1_5_en( T757 ),
       .io_VwirePorts_2_1_5_out( VwireModule_io_VwirePorts_2_1_5_out ),
       .io_VwirePorts_2_1_4_in( ArrayRowModule_2_io_V_wire_out_20 ),
       .io_VwirePorts_2_1_4_en( T756 ),
       .io_VwirePorts_2_1_4_out( VwireModule_io_VwirePorts_2_1_4_out ),
       .io_VwirePorts_2_1_3_in( ArrayRowModule_2_io_V_wire_out_19 ),
       .io_VwirePorts_2_1_3_en( T755 ),
       .io_VwirePorts_2_1_3_out( VwireModule_io_VwirePorts_2_1_3_out ),
       .io_VwirePorts_2_1_2_in( ArrayRowModule_2_io_V_wire_out_18 ),
       .io_VwirePorts_2_1_2_en( T754 ),
       .io_VwirePorts_2_1_2_out( VwireModule_io_VwirePorts_2_1_2_out ),
       .io_VwirePorts_2_1_1_in( ArrayRowModule_2_io_V_wire_out_17 ),
       .io_VwirePorts_2_1_1_en( T753 ),
       .io_VwirePorts_2_1_1_out( VwireModule_io_VwirePorts_2_1_1_out ),
       .io_VwirePorts_2_1_0_in( ArrayRowModule_2_io_V_wire_out_16 ),
       .io_VwirePorts_2_1_0_en( T752 ),
       .io_VwirePorts_2_1_0_out( VwireModule_io_VwirePorts_2_1_0_out ),
       .io_VwirePorts_2_0_15_in( ArrayRowModule_2_io_V_wire_out_15 ),
       .io_VwirePorts_2_0_15_en( T751 ),
       .io_VwirePorts_2_0_15_out( VwireModule_io_VwirePorts_2_0_15_out ),
       .io_VwirePorts_2_0_14_in( ArrayRowModule_2_io_V_wire_out_14 ),
       .io_VwirePorts_2_0_14_en( T750 ),
       .io_VwirePorts_2_0_14_out( VwireModule_io_VwirePorts_2_0_14_out ),
       .io_VwirePorts_2_0_13_in( ArrayRowModule_2_io_V_wire_out_13 ),
       .io_VwirePorts_2_0_13_en( T749 ),
       .io_VwirePorts_2_0_13_out( VwireModule_io_VwirePorts_2_0_13_out ),
       .io_VwirePorts_2_0_12_in( ArrayRowModule_2_io_V_wire_out_12 ),
       .io_VwirePorts_2_0_12_en( T748 ),
       .io_VwirePorts_2_0_12_out( VwireModule_io_VwirePorts_2_0_12_out ),
       .io_VwirePorts_2_0_11_in( ArrayRowModule_2_io_V_wire_out_11 ),
       .io_VwirePorts_2_0_11_en( T747 ),
       .io_VwirePorts_2_0_11_out( VwireModule_io_VwirePorts_2_0_11_out ),
       .io_VwirePorts_2_0_10_in( ArrayRowModule_2_io_V_wire_out_10 ),
       .io_VwirePorts_2_0_10_en( T746 ),
       .io_VwirePorts_2_0_10_out( VwireModule_io_VwirePorts_2_0_10_out ),
       .io_VwirePorts_2_0_9_in( ArrayRowModule_2_io_V_wire_out_9 ),
       .io_VwirePorts_2_0_9_en( T745 ),
       .io_VwirePorts_2_0_9_out( VwireModule_io_VwirePorts_2_0_9_out ),
       .io_VwirePorts_2_0_8_in( ArrayRowModule_2_io_V_wire_out_8 ),
       .io_VwirePorts_2_0_8_en( T744 ),
       .io_VwirePorts_2_0_8_out( VwireModule_io_VwirePorts_2_0_8_out ),
       .io_VwirePorts_2_0_7_in( ArrayRowModule_2_io_V_wire_out_7 ),
       .io_VwirePorts_2_0_7_en( T743 ),
       .io_VwirePorts_2_0_7_out( VwireModule_io_VwirePorts_2_0_7_out ),
       .io_VwirePorts_2_0_6_in( ArrayRowModule_2_io_V_wire_out_6 ),
       .io_VwirePorts_2_0_6_en( T742 ),
       .io_VwirePorts_2_0_6_out( VwireModule_io_VwirePorts_2_0_6_out ),
       .io_VwirePorts_2_0_5_in( ArrayRowModule_2_io_V_wire_out_5 ),
       .io_VwirePorts_2_0_5_en( T741 ),
       .io_VwirePorts_2_0_5_out( VwireModule_io_VwirePorts_2_0_5_out ),
       .io_VwirePorts_2_0_4_in( ArrayRowModule_2_io_V_wire_out_4 ),
       .io_VwirePorts_2_0_4_en( T740 ),
       .io_VwirePorts_2_0_4_out( VwireModule_io_VwirePorts_2_0_4_out ),
       .io_VwirePorts_2_0_3_in( ArrayRowModule_2_io_V_wire_out_3 ),
       .io_VwirePorts_2_0_3_en( T739 ),
       .io_VwirePorts_2_0_3_out( VwireModule_io_VwirePorts_2_0_3_out ),
       .io_VwirePorts_2_0_2_in( ArrayRowModule_2_io_V_wire_out_2 ),
       .io_VwirePorts_2_0_2_en( T738 ),
       .io_VwirePorts_2_0_2_out( VwireModule_io_VwirePorts_2_0_2_out ),
       .io_VwirePorts_2_0_1_in( ArrayRowModule_2_io_V_wire_out_1 ),
       .io_VwirePorts_2_0_1_en( T737 ),
       .io_VwirePorts_2_0_1_out( VwireModule_io_VwirePorts_2_0_1_out ),
       .io_VwirePorts_2_0_0_in( ArrayRowModule_2_io_V_wire_out_0 ),
       .io_VwirePorts_2_0_0_en( T736 ),
       .io_VwirePorts_2_0_0_out( VwireModule_io_VwirePorts_2_0_0_out ),
       .io_VwirePorts_1_22_15_in( ArrayRowModule_1_io_V_wire_out_367 ),
       .io_VwirePorts_1_22_15_en( T735 ),
       .io_VwirePorts_1_22_15_out( VwireModule_io_VwirePorts_1_22_15_out ),
       .io_VwirePorts_1_22_14_in( ArrayRowModule_1_io_V_wire_out_366 ),
       .io_VwirePorts_1_22_14_en( T734 ),
       .io_VwirePorts_1_22_14_out( VwireModule_io_VwirePorts_1_22_14_out ),
       .io_VwirePorts_1_22_13_in( ArrayRowModule_1_io_V_wire_out_365 ),
       .io_VwirePorts_1_22_13_en( T733 ),
       .io_VwirePorts_1_22_13_out( VwireModule_io_VwirePorts_1_22_13_out ),
       .io_VwirePorts_1_22_12_in( ArrayRowModule_1_io_V_wire_out_364 ),
       .io_VwirePorts_1_22_12_en( T732 ),
       .io_VwirePorts_1_22_12_out( VwireModule_io_VwirePorts_1_22_12_out ),
       .io_VwirePorts_1_22_11_in( ArrayRowModule_1_io_V_wire_out_363 ),
       .io_VwirePorts_1_22_11_en( T731 ),
       .io_VwirePorts_1_22_11_out( VwireModule_io_VwirePorts_1_22_11_out ),
       .io_VwirePorts_1_22_10_in( ArrayRowModule_1_io_V_wire_out_362 ),
       .io_VwirePorts_1_22_10_en( T730 ),
       .io_VwirePorts_1_22_10_out( VwireModule_io_VwirePorts_1_22_10_out ),
       .io_VwirePorts_1_22_9_in( ArrayRowModule_1_io_V_wire_out_361 ),
       .io_VwirePorts_1_22_9_en( T729 ),
       .io_VwirePorts_1_22_9_out( VwireModule_io_VwirePorts_1_22_9_out ),
       .io_VwirePorts_1_22_8_in( ArrayRowModule_1_io_V_wire_out_360 ),
       .io_VwirePorts_1_22_8_en( T728 ),
       .io_VwirePorts_1_22_8_out( VwireModule_io_VwirePorts_1_22_8_out ),
       .io_VwirePorts_1_22_7_in( ArrayRowModule_1_io_V_wire_out_359 ),
       .io_VwirePorts_1_22_7_en( T727 ),
       .io_VwirePorts_1_22_7_out( VwireModule_io_VwirePorts_1_22_7_out ),
       .io_VwirePorts_1_22_6_in( ArrayRowModule_1_io_V_wire_out_358 ),
       .io_VwirePorts_1_22_6_en( T726 ),
       .io_VwirePorts_1_22_6_out( VwireModule_io_VwirePorts_1_22_6_out ),
       .io_VwirePorts_1_22_5_in( ArrayRowModule_1_io_V_wire_out_357 ),
       .io_VwirePorts_1_22_5_en( T725 ),
       .io_VwirePorts_1_22_5_out( VwireModule_io_VwirePorts_1_22_5_out ),
       .io_VwirePorts_1_22_4_in( ArrayRowModule_1_io_V_wire_out_356 ),
       .io_VwirePorts_1_22_4_en( T724 ),
       .io_VwirePorts_1_22_4_out( VwireModule_io_VwirePorts_1_22_4_out ),
       .io_VwirePorts_1_22_3_in( ArrayRowModule_1_io_V_wire_out_355 ),
       .io_VwirePorts_1_22_3_en( T723 ),
       .io_VwirePorts_1_22_3_out( VwireModule_io_VwirePorts_1_22_3_out ),
       .io_VwirePorts_1_22_2_in( ArrayRowModule_1_io_V_wire_out_354 ),
       .io_VwirePorts_1_22_2_en( T722 ),
       .io_VwirePorts_1_22_2_out( VwireModule_io_VwirePorts_1_22_2_out ),
       .io_VwirePorts_1_22_1_in( ArrayRowModule_1_io_V_wire_out_353 ),
       .io_VwirePorts_1_22_1_en( T721 ),
       .io_VwirePorts_1_22_1_out( VwireModule_io_VwirePorts_1_22_1_out ),
       .io_VwirePorts_1_22_0_in( ArrayRowModule_1_io_V_wire_out_352 ),
       .io_VwirePorts_1_22_0_en( T720 ),
       .io_VwirePorts_1_22_0_out( VwireModule_io_VwirePorts_1_22_0_out ),
       .io_VwirePorts_1_21_15_in( ArrayRowModule_1_io_V_wire_out_351 ),
       .io_VwirePorts_1_21_15_en( T719 ),
       .io_VwirePorts_1_21_15_out( VwireModule_io_VwirePorts_1_21_15_out ),
       .io_VwirePorts_1_21_14_in( ArrayRowModule_1_io_V_wire_out_350 ),
       .io_VwirePorts_1_21_14_en( T718 ),
       .io_VwirePorts_1_21_14_out( VwireModule_io_VwirePorts_1_21_14_out ),
       .io_VwirePorts_1_21_13_in( ArrayRowModule_1_io_V_wire_out_349 ),
       .io_VwirePorts_1_21_13_en( T717 ),
       .io_VwirePorts_1_21_13_out( VwireModule_io_VwirePorts_1_21_13_out ),
       .io_VwirePorts_1_21_12_in( ArrayRowModule_1_io_V_wire_out_348 ),
       .io_VwirePorts_1_21_12_en( T716 ),
       .io_VwirePorts_1_21_12_out( VwireModule_io_VwirePorts_1_21_12_out ),
       .io_VwirePorts_1_21_11_in( ArrayRowModule_1_io_V_wire_out_347 ),
       .io_VwirePorts_1_21_11_en( T715 ),
       .io_VwirePorts_1_21_11_out( VwireModule_io_VwirePorts_1_21_11_out ),
       .io_VwirePorts_1_21_10_in( ArrayRowModule_1_io_V_wire_out_346 ),
       .io_VwirePorts_1_21_10_en( T714 ),
       .io_VwirePorts_1_21_10_out( VwireModule_io_VwirePorts_1_21_10_out ),
       .io_VwirePorts_1_21_9_in( ArrayRowModule_1_io_V_wire_out_345 ),
       .io_VwirePorts_1_21_9_en( T713 ),
       .io_VwirePorts_1_21_9_out( VwireModule_io_VwirePorts_1_21_9_out ),
       .io_VwirePorts_1_21_8_in( ArrayRowModule_1_io_V_wire_out_344 ),
       .io_VwirePorts_1_21_8_en( T712 ),
       .io_VwirePorts_1_21_8_out( VwireModule_io_VwirePorts_1_21_8_out ),
       .io_VwirePorts_1_21_7_in( ArrayRowModule_1_io_V_wire_out_343 ),
       .io_VwirePorts_1_21_7_en( T711 ),
       .io_VwirePorts_1_21_7_out( VwireModule_io_VwirePorts_1_21_7_out ),
       .io_VwirePorts_1_21_6_in( ArrayRowModule_1_io_V_wire_out_342 ),
       .io_VwirePorts_1_21_6_en( T710 ),
       .io_VwirePorts_1_21_6_out( VwireModule_io_VwirePorts_1_21_6_out ),
       .io_VwirePorts_1_21_5_in( ArrayRowModule_1_io_V_wire_out_341 ),
       .io_VwirePorts_1_21_5_en( T709 ),
       .io_VwirePorts_1_21_5_out( VwireModule_io_VwirePorts_1_21_5_out ),
       .io_VwirePorts_1_21_4_in( ArrayRowModule_1_io_V_wire_out_340 ),
       .io_VwirePorts_1_21_4_en( T708 ),
       .io_VwirePorts_1_21_4_out( VwireModule_io_VwirePorts_1_21_4_out ),
       .io_VwirePorts_1_21_3_in( ArrayRowModule_1_io_V_wire_out_339 ),
       .io_VwirePorts_1_21_3_en( T707 ),
       .io_VwirePorts_1_21_3_out( VwireModule_io_VwirePorts_1_21_3_out ),
       .io_VwirePorts_1_21_2_in( ArrayRowModule_1_io_V_wire_out_338 ),
       .io_VwirePorts_1_21_2_en( T706 ),
       .io_VwirePorts_1_21_2_out( VwireModule_io_VwirePorts_1_21_2_out ),
       .io_VwirePorts_1_21_1_in( ArrayRowModule_1_io_V_wire_out_337 ),
       .io_VwirePorts_1_21_1_en( T705 ),
       .io_VwirePorts_1_21_1_out( VwireModule_io_VwirePorts_1_21_1_out ),
       .io_VwirePorts_1_21_0_in( ArrayRowModule_1_io_V_wire_out_336 ),
       .io_VwirePorts_1_21_0_en( T704 ),
       .io_VwirePorts_1_21_0_out( VwireModule_io_VwirePorts_1_21_0_out ),
       .io_VwirePorts_1_20_15_in( ArrayRowModule_1_io_V_wire_out_335 ),
       .io_VwirePorts_1_20_15_en( T703 ),
       .io_VwirePorts_1_20_15_out( VwireModule_io_VwirePorts_1_20_15_out ),
       .io_VwirePorts_1_20_14_in( ArrayRowModule_1_io_V_wire_out_334 ),
       .io_VwirePorts_1_20_14_en( T702 ),
       .io_VwirePorts_1_20_14_out( VwireModule_io_VwirePorts_1_20_14_out ),
       .io_VwirePorts_1_20_13_in( ArrayRowModule_1_io_V_wire_out_333 ),
       .io_VwirePorts_1_20_13_en( T701 ),
       .io_VwirePorts_1_20_13_out( VwireModule_io_VwirePorts_1_20_13_out ),
       .io_VwirePorts_1_20_12_in( ArrayRowModule_1_io_V_wire_out_332 ),
       .io_VwirePorts_1_20_12_en( T700 ),
       .io_VwirePorts_1_20_12_out( VwireModule_io_VwirePorts_1_20_12_out ),
       .io_VwirePorts_1_20_11_in( ArrayRowModule_1_io_V_wire_out_331 ),
       .io_VwirePorts_1_20_11_en( T699 ),
       .io_VwirePorts_1_20_11_out( VwireModule_io_VwirePorts_1_20_11_out ),
       .io_VwirePorts_1_20_10_in( ArrayRowModule_1_io_V_wire_out_330 ),
       .io_VwirePorts_1_20_10_en( T698 ),
       .io_VwirePorts_1_20_10_out( VwireModule_io_VwirePorts_1_20_10_out ),
       .io_VwirePorts_1_20_9_in( ArrayRowModule_1_io_V_wire_out_329 ),
       .io_VwirePorts_1_20_9_en( T697 ),
       .io_VwirePorts_1_20_9_out( VwireModule_io_VwirePorts_1_20_9_out ),
       .io_VwirePorts_1_20_8_in( ArrayRowModule_1_io_V_wire_out_328 ),
       .io_VwirePorts_1_20_8_en( T696 ),
       .io_VwirePorts_1_20_8_out( VwireModule_io_VwirePorts_1_20_8_out ),
       .io_VwirePorts_1_20_7_in( ArrayRowModule_1_io_V_wire_out_327 ),
       .io_VwirePorts_1_20_7_en( T695 ),
       .io_VwirePorts_1_20_7_out( VwireModule_io_VwirePorts_1_20_7_out ),
       .io_VwirePorts_1_20_6_in( ArrayRowModule_1_io_V_wire_out_326 ),
       .io_VwirePorts_1_20_6_en( T694 ),
       .io_VwirePorts_1_20_6_out( VwireModule_io_VwirePorts_1_20_6_out ),
       .io_VwirePorts_1_20_5_in( ArrayRowModule_1_io_V_wire_out_325 ),
       .io_VwirePorts_1_20_5_en( T693 ),
       .io_VwirePorts_1_20_5_out( VwireModule_io_VwirePorts_1_20_5_out ),
       .io_VwirePorts_1_20_4_in( ArrayRowModule_1_io_V_wire_out_324 ),
       .io_VwirePorts_1_20_4_en( T692 ),
       .io_VwirePorts_1_20_4_out( VwireModule_io_VwirePorts_1_20_4_out ),
       .io_VwirePorts_1_20_3_in( ArrayRowModule_1_io_V_wire_out_323 ),
       .io_VwirePorts_1_20_3_en( T691 ),
       .io_VwirePorts_1_20_3_out( VwireModule_io_VwirePorts_1_20_3_out ),
       .io_VwirePorts_1_20_2_in( ArrayRowModule_1_io_V_wire_out_322 ),
       .io_VwirePorts_1_20_2_en( T690 ),
       .io_VwirePorts_1_20_2_out( VwireModule_io_VwirePorts_1_20_2_out ),
       .io_VwirePorts_1_20_1_in( ArrayRowModule_1_io_V_wire_out_321 ),
       .io_VwirePorts_1_20_1_en( T689 ),
       .io_VwirePorts_1_20_1_out( VwireModule_io_VwirePorts_1_20_1_out ),
       .io_VwirePorts_1_20_0_in( ArrayRowModule_1_io_V_wire_out_320 ),
       .io_VwirePorts_1_20_0_en( T688 ),
       .io_VwirePorts_1_20_0_out( VwireModule_io_VwirePorts_1_20_0_out ),
       .io_VwirePorts_1_19_15_in( ArrayRowModule_1_io_V_wire_out_319 ),
       .io_VwirePorts_1_19_15_en( T687 ),
       .io_VwirePorts_1_19_15_out( VwireModule_io_VwirePorts_1_19_15_out ),
       .io_VwirePorts_1_19_14_in( ArrayRowModule_1_io_V_wire_out_318 ),
       .io_VwirePorts_1_19_14_en( T686 ),
       .io_VwirePorts_1_19_14_out( VwireModule_io_VwirePorts_1_19_14_out ),
       .io_VwirePorts_1_19_13_in( ArrayRowModule_1_io_V_wire_out_317 ),
       .io_VwirePorts_1_19_13_en( T685 ),
       .io_VwirePorts_1_19_13_out( VwireModule_io_VwirePorts_1_19_13_out ),
       .io_VwirePorts_1_19_12_in( ArrayRowModule_1_io_V_wire_out_316 ),
       .io_VwirePorts_1_19_12_en( T684 ),
       .io_VwirePorts_1_19_12_out( VwireModule_io_VwirePorts_1_19_12_out ),
       .io_VwirePorts_1_19_11_in( ArrayRowModule_1_io_V_wire_out_315 ),
       .io_VwirePorts_1_19_11_en( T683 ),
       .io_VwirePorts_1_19_11_out( VwireModule_io_VwirePorts_1_19_11_out ),
       .io_VwirePorts_1_19_10_in( ArrayRowModule_1_io_V_wire_out_314 ),
       .io_VwirePorts_1_19_10_en( T682 ),
       .io_VwirePorts_1_19_10_out( VwireModule_io_VwirePorts_1_19_10_out ),
       .io_VwirePorts_1_19_9_in( ArrayRowModule_1_io_V_wire_out_313 ),
       .io_VwirePorts_1_19_9_en( T681 ),
       .io_VwirePorts_1_19_9_out( VwireModule_io_VwirePorts_1_19_9_out ),
       .io_VwirePorts_1_19_8_in( ArrayRowModule_1_io_V_wire_out_312 ),
       .io_VwirePorts_1_19_8_en( T680 ),
       .io_VwirePorts_1_19_8_out( VwireModule_io_VwirePorts_1_19_8_out ),
       .io_VwirePorts_1_19_7_in( ArrayRowModule_1_io_V_wire_out_311 ),
       .io_VwirePorts_1_19_7_en( T679 ),
       .io_VwirePorts_1_19_7_out( VwireModule_io_VwirePorts_1_19_7_out ),
       .io_VwirePorts_1_19_6_in( ArrayRowModule_1_io_V_wire_out_310 ),
       .io_VwirePorts_1_19_6_en( T678 ),
       .io_VwirePorts_1_19_6_out( VwireModule_io_VwirePorts_1_19_6_out ),
       .io_VwirePorts_1_19_5_in( ArrayRowModule_1_io_V_wire_out_309 ),
       .io_VwirePorts_1_19_5_en( T677 ),
       .io_VwirePorts_1_19_5_out( VwireModule_io_VwirePorts_1_19_5_out ),
       .io_VwirePorts_1_19_4_in( ArrayRowModule_1_io_V_wire_out_308 ),
       .io_VwirePorts_1_19_4_en( T676 ),
       .io_VwirePorts_1_19_4_out( VwireModule_io_VwirePorts_1_19_4_out ),
       .io_VwirePorts_1_19_3_in( ArrayRowModule_1_io_V_wire_out_307 ),
       .io_VwirePorts_1_19_3_en( T675 ),
       .io_VwirePorts_1_19_3_out( VwireModule_io_VwirePorts_1_19_3_out ),
       .io_VwirePorts_1_19_2_in( ArrayRowModule_1_io_V_wire_out_306 ),
       .io_VwirePorts_1_19_2_en( T674 ),
       .io_VwirePorts_1_19_2_out( VwireModule_io_VwirePorts_1_19_2_out ),
       .io_VwirePorts_1_19_1_in( ArrayRowModule_1_io_V_wire_out_305 ),
       .io_VwirePorts_1_19_1_en( T673 ),
       .io_VwirePorts_1_19_1_out( VwireModule_io_VwirePorts_1_19_1_out ),
       .io_VwirePorts_1_19_0_in( ArrayRowModule_1_io_V_wire_out_304 ),
       .io_VwirePorts_1_19_0_en( T672 ),
       .io_VwirePorts_1_19_0_out( VwireModule_io_VwirePorts_1_19_0_out ),
       .io_VwirePorts_1_18_15_in( ArrayRowModule_1_io_V_wire_out_303 ),
       .io_VwirePorts_1_18_15_en( T671 ),
       .io_VwirePorts_1_18_15_out( VwireModule_io_VwirePorts_1_18_15_out ),
       .io_VwirePorts_1_18_14_in( ArrayRowModule_1_io_V_wire_out_302 ),
       .io_VwirePorts_1_18_14_en( T670 ),
       .io_VwirePorts_1_18_14_out( VwireModule_io_VwirePorts_1_18_14_out ),
       .io_VwirePorts_1_18_13_in( ArrayRowModule_1_io_V_wire_out_301 ),
       .io_VwirePorts_1_18_13_en( T669 ),
       .io_VwirePorts_1_18_13_out( VwireModule_io_VwirePorts_1_18_13_out ),
       .io_VwirePorts_1_18_12_in( ArrayRowModule_1_io_V_wire_out_300 ),
       .io_VwirePorts_1_18_12_en( T668 ),
       .io_VwirePorts_1_18_12_out( VwireModule_io_VwirePorts_1_18_12_out ),
       .io_VwirePorts_1_18_11_in( ArrayRowModule_1_io_V_wire_out_299 ),
       .io_VwirePorts_1_18_11_en( T667 ),
       .io_VwirePorts_1_18_11_out( VwireModule_io_VwirePorts_1_18_11_out ),
       .io_VwirePorts_1_18_10_in( ArrayRowModule_1_io_V_wire_out_298 ),
       .io_VwirePorts_1_18_10_en( T666 ),
       .io_VwirePorts_1_18_10_out( VwireModule_io_VwirePorts_1_18_10_out ),
       .io_VwirePorts_1_18_9_in( ArrayRowModule_1_io_V_wire_out_297 ),
       .io_VwirePorts_1_18_9_en( T665 ),
       .io_VwirePorts_1_18_9_out( VwireModule_io_VwirePorts_1_18_9_out ),
       .io_VwirePorts_1_18_8_in( ArrayRowModule_1_io_V_wire_out_296 ),
       .io_VwirePorts_1_18_8_en( T664 ),
       .io_VwirePorts_1_18_8_out( VwireModule_io_VwirePorts_1_18_8_out ),
       .io_VwirePorts_1_18_7_in( ArrayRowModule_1_io_V_wire_out_295 ),
       .io_VwirePorts_1_18_7_en( T663 ),
       .io_VwirePorts_1_18_7_out( VwireModule_io_VwirePorts_1_18_7_out ),
       .io_VwirePorts_1_18_6_in( ArrayRowModule_1_io_V_wire_out_294 ),
       .io_VwirePorts_1_18_6_en( T662 ),
       .io_VwirePorts_1_18_6_out( VwireModule_io_VwirePorts_1_18_6_out ),
       .io_VwirePorts_1_18_5_in( ArrayRowModule_1_io_V_wire_out_293 ),
       .io_VwirePorts_1_18_5_en( T661 ),
       .io_VwirePorts_1_18_5_out( VwireModule_io_VwirePorts_1_18_5_out ),
       .io_VwirePorts_1_18_4_in( ArrayRowModule_1_io_V_wire_out_292 ),
       .io_VwirePorts_1_18_4_en( T660 ),
       .io_VwirePorts_1_18_4_out( VwireModule_io_VwirePorts_1_18_4_out ),
       .io_VwirePorts_1_18_3_in( ArrayRowModule_1_io_V_wire_out_291 ),
       .io_VwirePorts_1_18_3_en( T659 ),
       .io_VwirePorts_1_18_3_out( VwireModule_io_VwirePorts_1_18_3_out ),
       .io_VwirePorts_1_18_2_in( ArrayRowModule_1_io_V_wire_out_290 ),
       .io_VwirePorts_1_18_2_en( T658 ),
       .io_VwirePorts_1_18_2_out( VwireModule_io_VwirePorts_1_18_2_out ),
       .io_VwirePorts_1_18_1_in( ArrayRowModule_1_io_V_wire_out_289 ),
       .io_VwirePorts_1_18_1_en( T657 ),
       .io_VwirePorts_1_18_1_out( VwireModule_io_VwirePorts_1_18_1_out ),
       .io_VwirePorts_1_18_0_in( ArrayRowModule_1_io_V_wire_out_288 ),
       .io_VwirePorts_1_18_0_en( T656 ),
       .io_VwirePorts_1_18_0_out( VwireModule_io_VwirePorts_1_18_0_out ),
       .io_VwirePorts_1_17_15_in( ArrayRowModule_1_io_V_wire_out_287 ),
       .io_VwirePorts_1_17_15_en( T655 ),
       .io_VwirePorts_1_17_15_out( VwireModule_io_VwirePorts_1_17_15_out ),
       .io_VwirePorts_1_17_14_in( ArrayRowModule_1_io_V_wire_out_286 ),
       .io_VwirePorts_1_17_14_en( T654 ),
       .io_VwirePorts_1_17_14_out( VwireModule_io_VwirePorts_1_17_14_out ),
       .io_VwirePorts_1_17_13_in( ArrayRowModule_1_io_V_wire_out_285 ),
       .io_VwirePorts_1_17_13_en( T653 ),
       .io_VwirePorts_1_17_13_out( VwireModule_io_VwirePorts_1_17_13_out ),
       .io_VwirePorts_1_17_12_in( ArrayRowModule_1_io_V_wire_out_284 ),
       .io_VwirePorts_1_17_12_en( T652 ),
       .io_VwirePorts_1_17_12_out( VwireModule_io_VwirePorts_1_17_12_out ),
       .io_VwirePorts_1_17_11_in( ArrayRowModule_1_io_V_wire_out_283 ),
       .io_VwirePorts_1_17_11_en( T651 ),
       .io_VwirePorts_1_17_11_out( VwireModule_io_VwirePorts_1_17_11_out ),
       .io_VwirePorts_1_17_10_in( ArrayRowModule_1_io_V_wire_out_282 ),
       .io_VwirePorts_1_17_10_en( T650 ),
       .io_VwirePorts_1_17_10_out( VwireModule_io_VwirePorts_1_17_10_out ),
       .io_VwirePorts_1_17_9_in( ArrayRowModule_1_io_V_wire_out_281 ),
       .io_VwirePorts_1_17_9_en( T649 ),
       .io_VwirePorts_1_17_9_out( VwireModule_io_VwirePorts_1_17_9_out ),
       .io_VwirePorts_1_17_8_in( ArrayRowModule_1_io_V_wire_out_280 ),
       .io_VwirePorts_1_17_8_en( T648 ),
       .io_VwirePorts_1_17_8_out( VwireModule_io_VwirePorts_1_17_8_out ),
       .io_VwirePorts_1_17_7_in( ArrayRowModule_1_io_V_wire_out_279 ),
       .io_VwirePorts_1_17_7_en( T647 ),
       .io_VwirePorts_1_17_7_out( VwireModule_io_VwirePorts_1_17_7_out ),
       .io_VwirePorts_1_17_6_in( ArrayRowModule_1_io_V_wire_out_278 ),
       .io_VwirePorts_1_17_6_en( T646 ),
       .io_VwirePorts_1_17_6_out( VwireModule_io_VwirePorts_1_17_6_out ),
       .io_VwirePorts_1_17_5_in( ArrayRowModule_1_io_V_wire_out_277 ),
       .io_VwirePorts_1_17_5_en( T645 ),
       .io_VwirePorts_1_17_5_out( VwireModule_io_VwirePorts_1_17_5_out ),
       .io_VwirePorts_1_17_4_in( ArrayRowModule_1_io_V_wire_out_276 ),
       .io_VwirePorts_1_17_4_en( T644 ),
       .io_VwirePorts_1_17_4_out( VwireModule_io_VwirePorts_1_17_4_out ),
       .io_VwirePorts_1_17_3_in( ArrayRowModule_1_io_V_wire_out_275 ),
       .io_VwirePorts_1_17_3_en( T643 ),
       .io_VwirePorts_1_17_3_out( VwireModule_io_VwirePorts_1_17_3_out ),
       .io_VwirePorts_1_17_2_in( ArrayRowModule_1_io_V_wire_out_274 ),
       .io_VwirePorts_1_17_2_en( T642 ),
       .io_VwirePorts_1_17_2_out( VwireModule_io_VwirePorts_1_17_2_out ),
       .io_VwirePorts_1_17_1_in( ArrayRowModule_1_io_V_wire_out_273 ),
       .io_VwirePorts_1_17_1_en( T641 ),
       .io_VwirePorts_1_17_1_out( VwireModule_io_VwirePorts_1_17_1_out ),
       .io_VwirePorts_1_17_0_in( ArrayRowModule_1_io_V_wire_out_272 ),
       .io_VwirePorts_1_17_0_en( T640 ),
       .io_VwirePorts_1_17_0_out( VwireModule_io_VwirePorts_1_17_0_out ),
       .io_VwirePorts_1_16_15_in( ArrayRowModule_1_io_V_wire_out_271 ),
       .io_VwirePorts_1_16_15_en( T639 ),
       .io_VwirePorts_1_16_15_out( VwireModule_io_VwirePorts_1_16_15_out ),
       .io_VwirePorts_1_16_14_in( ArrayRowModule_1_io_V_wire_out_270 ),
       .io_VwirePorts_1_16_14_en( T638 ),
       .io_VwirePorts_1_16_14_out( VwireModule_io_VwirePorts_1_16_14_out ),
       .io_VwirePorts_1_16_13_in( ArrayRowModule_1_io_V_wire_out_269 ),
       .io_VwirePorts_1_16_13_en( T637 ),
       .io_VwirePorts_1_16_13_out( VwireModule_io_VwirePorts_1_16_13_out ),
       .io_VwirePorts_1_16_12_in( ArrayRowModule_1_io_V_wire_out_268 ),
       .io_VwirePorts_1_16_12_en( T636 ),
       .io_VwirePorts_1_16_12_out( VwireModule_io_VwirePorts_1_16_12_out ),
       .io_VwirePorts_1_16_11_in( ArrayRowModule_1_io_V_wire_out_267 ),
       .io_VwirePorts_1_16_11_en( T635 ),
       .io_VwirePorts_1_16_11_out( VwireModule_io_VwirePorts_1_16_11_out ),
       .io_VwirePorts_1_16_10_in( ArrayRowModule_1_io_V_wire_out_266 ),
       .io_VwirePorts_1_16_10_en( T634 ),
       .io_VwirePorts_1_16_10_out( VwireModule_io_VwirePorts_1_16_10_out ),
       .io_VwirePorts_1_16_9_in( ArrayRowModule_1_io_V_wire_out_265 ),
       .io_VwirePorts_1_16_9_en( T633 ),
       .io_VwirePorts_1_16_9_out( VwireModule_io_VwirePorts_1_16_9_out ),
       .io_VwirePorts_1_16_8_in( ArrayRowModule_1_io_V_wire_out_264 ),
       .io_VwirePorts_1_16_8_en( T632 ),
       .io_VwirePorts_1_16_8_out( VwireModule_io_VwirePorts_1_16_8_out ),
       .io_VwirePorts_1_16_7_in( ArrayRowModule_1_io_V_wire_out_263 ),
       .io_VwirePorts_1_16_7_en( T631 ),
       .io_VwirePorts_1_16_7_out( VwireModule_io_VwirePorts_1_16_7_out ),
       .io_VwirePorts_1_16_6_in( ArrayRowModule_1_io_V_wire_out_262 ),
       .io_VwirePorts_1_16_6_en( T630 ),
       .io_VwirePorts_1_16_6_out( VwireModule_io_VwirePorts_1_16_6_out ),
       .io_VwirePorts_1_16_5_in( ArrayRowModule_1_io_V_wire_out_261 ),
       .io_VwirePorts_1_16_5_en( T629 ),
       .io_VwirePorts_1_16_5_out( VwireModule_io_VwirePorts_1_16_5_out ),
       .io_VwirePorts_1_16_4_in( ArrayRowModule_1_io_V_wire_out_260 ),
       .io_VwirePorts_1_16_4_en( T628 ),
       .io_VwirePorts_1_16_4_out( VwireModule_io_VwirePorts_1_16_4_out ),
       .io_VwirePorts_1_16_3_in( ArrayRowModule_1_io_V_wire_out_259 ),
       .io_VwirePorts_1_16_3_en( T627 ),
       .io_VwirePorts_1_16_3_out( VwireModule_io_VwirePorts_1_16_3_out ),
       .io_VwirePorts_1_16_2_in( ArrayRowModule_1_io_V_wire_out_258 ),
       .io_VwirePorts_1_16_2_en( T626 ),
       .io_VwirePorts_1_16_2_out( VwireModule_io_VwirePorts_1_16_2_out ),
       .io_VwirePorts_1_16_1_in( ArrayRowModule_1_io_V_wire_out_257 ),
       .io_VwirePorts_1_16_1_en( T625 ),
       .io_VwirePorts_1_16_1_out( VwireModule_io_VwirePorts_1_16_1_out ),
       .io_VwirePorts_1_16_0_in( ArrayRowModule_1_io_V_wire_out_256 ),
       .io_VwirePorts_1_16_0_en( T624 ),
       .io_VwirePorts_1_16_0_out( VwireModule_io_VwirePorts_1_16_0_out ),
       .io_VwirePorts_1_15_15_in( ArrayRowModule_1_io_V_wire_out_255 ),
       .io_VwirePorts_1_15_15_en( T623 ),
       .io_VwirePorts_1_15_15_out( VwireModule_io_VwirePorts_1_15_15_out ),
       .io_VwirePorts_1_15_14_in( ArrayRowModule_1_io_V_wire_out_254 ),
       .io_VwirePorts_1_15_14_en( T622 ),
       .io_VwirePorts_1_15_14_out( VwireModule_io_VwirePorts_1_15_14_out ),
       .io_VwirePorts_1_15_13_in( ArrayRowModule_1_io_V_wire_out_253 ),
       .io_VwirePorts_1_15_13_en( T621 ),
       .io_VwirePorts_1_15_13_out( VwireModule_io_VwirePorts_1_15_13_out ),
       .io_VwirePorts_1_15_12_in( ArrayRowModule_1_io_V_wire_out_252 ),
       .io_VwirePorts_1_15_12_en( T620 ),
       .io_VwirePorts_1_15_12_out( VwireModule_io_VwirePorts_1_15_12_out ),
       .io_VwirePorts_1_15_11_in( ArrayRowModule_1_io_V_wire_out_251 ),
       .io_VwirePorts_1_15_11_en( T619 ),
       .io_VwirePorts_1_15_11_out( VwireModule_io_VwirePorts_1_15_11_out ),
       .io_VwirePorts_1_15_10_in( ArrayRowModule_1_io_V_wire_out_250 ),
       .io_VwirePorts_1_15_10_en( T618 ),
       .io_VwirePorts_1_15_10_out( VwireModule_io_VwirePorts_1_15_10_out ),
       .io_VwirePorts_1_15_9_in( ArrayRowModule_1_io_V_wire_out_249 ),
       .io_VwirePorts_1_15_9_en( T617 ),
       .io_VwirePorts_1_15_9_out( VwireModule_io_VwirePorts_1_15_9_out ),
       .io_VwirePorts_1_15_8_in( ArrayRowModule_1_io_V_wire_out_248 ),
       .io_VwirePorts_1_15_8_en( T616 ),
       .io_VwirePorts_1_15_8_out( VwireModule_io_VwirePorts_1_15_8_out ),
       .io_VwirePorts_1_15_7_in( ArrayRowModule_1_io_V_wire_out_247 ),
       .io_VwirePorts_1_15_7_en( T615 ),
       .io_VwirePorts_1_15_7_out( VwireModule_io_VwirePorts_1_15_7_out ),
       .io_VwirePorts_1_15_6_in( ArrayRowModule_1_io_V_wire_out_246 ),
       .io_VwirePorts_1_15_6_en( T614 ),
       .io_VwirePorts_1_15_6_out( VwireModule_io_VwirePorts_1_15_6_out ),
       .io_VwirePorts_1_15_5_in( ArrayRowModule_1_io_V_wire_out_245 ),
       .io_VwirePorts_1_15_5_en( T613 ),
       .io_VwirePorts_1_15_5_out( VwireModule_io_VwirePorts_1_15_5_out ),
       .io_VwirePorts_1_15_4_in( ArrayRowModule_1_io_V_wire_out_244 ),
       .io_VwirePorts_1_15_4_en( T612 ),
       .io_VwirePorts_1_15_4_out( VwireModule_io_VwirePorts_1_15_4_out ),
       .io_VwirePorts_1_15_3_in( ArrayRowModule_1_io_V_wire_out_243 ),
       .io_VwirePorts_1_15_3_en( T611 ),
       .io_VwirePorts_1_15_3_out( VwireModule_io_VwirePorts_1_15_3_out ),
       .io_VwirePorts_1_15_2_in( ArrayRowModule_1_io_V_wire_out_242 ),
       .io_VwirePorts_1_15_2_en( T610 ),
       .io_VwirePorts_1_15_2_out( VwireModule_io_VwirePorts_1_15_2_out ),
       .io_VwirePorts_1_15_1_in( ArrayRowModule_1_io_V_wire_out_241 ),
       .io_VwirePorts_1_15_1_en( T609 ),
       .io_VwirePorts_1_15_1_out( VwireModule_io_VwirePorts_1_15_1_out ),
       .io_VwirePorts_1_15_0_in( ArrayRowModule_1_io_V_wire_out_240 ),
       .io_VwirePorts_1_15_0_en( T608 ),
       .io_VwirePorts_1_15_0_out( VwireModule_io_VwirePorts_1_15_0_out ),
       .io_VwirePorts_1_14_15_in( ArrayRowModule_1_io_V_wire_out_239 ),
       .io_VwirePorts_1_14_15_en( T607 ),
       .io_VwirePorts_1_14_15_out( VwireModule_io_VwirePorts_1_14_15_out ),
       .io_VwirePorts_1_14_14_in( ArrayRowModule_1_io_V_wire_out_238 ),
       .io_VwirePorts_1_14_14_en( T606 ),
       .io_VwirePorts_1_14_14_out( VwireModule_io_VwirePorts_1_14_14_out ),
       .io_VwirePorts_1_14_13_in( ArrayRowModule_1_io_V_wire_out_237 ),
       .io_VwirePorts_1_14_13_en( T605 ),
       .io_VwirePorts_1_14_13_out( VwireModule_io_VwirePorts_1_14_13_out ),
       .io_VwirePorts_1_14_12_in( ArrayRowModule_1_io_V_wire_out_236 ),
       .io_VwirePorts_1_14_12_en( T604 ),
       .io_VwirePorts_1_14_12_out( VwireModule_io_VwirePorts_1_14_12_out ),
       .io_VwirePorts_1_14_11_in( ArrayRowModule_1_io_V_wire_out_235 ),
       .io_VwirePorts_1_14_11_en( T603 ),
       .io_VwirePorts_1_14_11_out( VwireModule_io_VwirePorts_1_14_11_out ),
       .io_VwirePorts_1_14_10_in( ArrayRowModule_1_io_V_wire_out_234 ),
       .io_VwirePorts_1_14_10_en( T602 ),
       .io_VwirePorts_1_14_10_out( VwireModule_io_VwirePorts_1_14_10_out ),
       .io_VwirePorts_1_14_9_in( ArrayRowModule_1_io_V_wire_out_233 ),
       .io_VwirePorts_1_14_9_en( T601 ),
       .io_VwirePorts_1_14_9_out( VwireModule_io_VwirePorts_1_14_9_out ),
       .io_VwirePorts_1_14_8_in( ArrayRowModule_1_io_V_wire_out_232 ),
       .io_VwirePorts_1_14_8_en( T600 ),
       .io_VwirePorts_1_14_8_out( VwireModule_io_VwirePorts_1_14_8_out ),
       .io_VwirePorts_1_14_7_in( ArrayRowModule_1_io_V_wire_out_231 ),
       .io_VwirePorts_1_14_7_en( T599 ),
       .io_VwirePorts_1_14_7_out( VwireModule_io_VwirePorts_1_14_7_out ),
       .io_VwirePorts_1_14_6_in( ArrayRowModule_1_io_V_wire_out_230 ),
       .io_VwirePorts_1_14_6_en( T598 ),
       .io_VwirePorts_1_14_6_out( VwireModule_io_VwirePorts_1_14_6_out ),
       .io_VwirePorts_1_14_5_in( ArrayRowModule_1_io_V_wire_out_229 ),
       .io_VwirePorts_1_14_5_en( T597 ),
       .io_VwirePorts_1_14_5_out( VwireModule_io_VwirePorts_1_14_5_out ),
       .io_VwirePorts_1_14_4_in( ArrayRowModule_1_io_V_wire_out_228 ),
       .io_VwirePorts_1_14_4_en( T596 ),
       .io_VwirePorts_1_14_4_out( VwireModule_io_VwirePorts_1_14_4_out ),
       .io_VwirePorts_1_14_3_in( ArrayRowModule_1_io_V_wire_out_227 ),
       .io_VwirePorts_1_14_3_en( T595 ),
       .io_VwirePorts_1_14_3_out( VwireModule_io_VwirePorts_1_14_3_out ),
       .io_VwirePorts_1_14_2_in( ArrayRowModule_1_io_V_wire_out_226 ),
       .io_VwirePorts_1_14_2_en( T594 ),
       .io_VwirePorts_1_14_2_out( VwireModule_io_VwirePorts_1_14_2_out ),
       .io_VwirePorts_1_14_1_in( ArrayRowModule_1_io_V_wire_out_225 ),
       .io_VwirePorts_1_14_1_en( T593 ),
       .io_VwirePorts_1_14_1_out( VwireModule_io_VwirePorts_1_14_1_out ),
       .io_VwirePorts_1_14_0_in( ArrayRowModule_1_io_V_wire_out_224 ),
       .io_VwirePorts_1_14_0_en( T592 ),
       .io_VwirePorts_1_14_0_out( VwireModule_io_VwirePorts_1_14_0_out ),
       .io_VwirePorts_1_13_15_in( ArrayRowModule_1_io_V_wire_out_223 ),
       .io_VwirePorts_1_13_15_en( T591 ),
       .io_VwirePorts_1_13_15_out( VwireModule_io_VwirePorts_1_13_15_out ),
       .io_VwirePorts_1_13_14_in( ArrayRowModule_1_io_V_wire_out_222 ),
       .io_VwirePorts_1_13_14_en( T590 ),
       .io_VwirePorts_1_13_14_out( VwireModule_io_VwirePorts_1_13_14_out ),
       .io_VwirePorts_1_13_13_in( ArrayRowModule_1_io_V_wire_out_221 ),
       .io_VwirePorts_1_13_13_en( T589 ),
       .io_VwirePorts_1_13_13_out( VwireModule_io_VwirePorts_1_13_13_out ),
       .io_VwirePorts_1_13_12_in( ArrayRowModule_1_io_V_wire_out_220 ),
       .io_VwirePorts_1_13_12_en( T588 ),
       .io_VwirePorts_1_13_12_out( VwireModule_io_VwirePorts_1_13_12_out ),
       .io_VwirePorts_1_13_11_in( ArrayRowModule_1_io_V_wire_out_219 ),
       .io_VwirePorts_1_13_11_en( T587 ),
       .io_VwirePorts_1_13_11_out( VwireModule_io_VwirePorts_1_13_11_out ),
       .io_VwirePorts_1_13_10_in( ArrayRowModule_1_io_V_wire_out_218 ),
       .io_VwirePorts_1_13_10_en( T586 ),
       .io_VwirePorts_1_13_10_out( VwireModule_io_VwirePorts_1_13_10_out ),
       .io_VwirePorts_1_13_9_in( ArrayRowModule_1_io_V_wire_out_217 ),
       .io_VwirePorts_1_13_9_en( T585 ),
       .io_VwirePorts_1_13_9_out( VwireModule_io_VwirePorts_1_13_9_out ),
       .io_VwirePorts_1_13_8_in( ArrayRowModule_1_io_V_wire_out_216 ),
       .io_VwirePorts_1_13_8_en( T584 ),
       .io_VwirePorts_1_13_8_out( VwireModule_io_VwirePorts_1_13_8_out ),
       .io_VwirePorts_1_13_7_in( ArrayRowModule_1_io_V_wire_out_215 ),
       .io_VwirePorts_1_13_7_en( T583 ),
       .io_VwirePorts_1_13_7_out( VwireModule_io_VwirePorts_1_13_7_out ),
       .io_VwirePorts_1_13_6_in( ArrayRowModule_1_io_V_wire_out_214 ),
       .io_VwirePorts_1_13_6_en( T582 ),
       .io_VwirePorts_1_13_6_out( VwireModule_io_VwirePorts_1_13_6_out ),
       .io_VwirePorts_1_13_5_in( ArrayRowModule_1_io_V_wire_out_213 ),
       .io_VwirePorts_1_13_5_en( T581 ),
       .io_VwirePorts_1_13_5_out( VwireModule_io_VwirePorts_1_13_5_out ),
       .io_VwirePorts_1_13_4_in( ArrayRowModule_1_io_V_wire_out_212 ),
       .io_VwirePorts_1_13_4_en( T580 ),
       .io_VwirePorts_1_13_4_out( VwireModule_io_VwirePorts_1_13_4_out ),
       .io_VwirePorts_1_13_3_in( ArrayRowModule_1_io_V_wire_out_211 ),
       .io_VwirePorts_1_13_3_en( T579 ),
       .io_VwirePorts_1_13_3_out( VwireModule_io_VwirePorts_1_13_3_out ),
       .io_VwirePorts_1_13_2_in( ArrayRowModule_1_io_V_wire_out_210 ),
       .io_VwirePorts_1_13_2_en( T578 ),
       .io_VwirePorts_1_13_2_out( VwireModule_io_VwirePorts_1_13_2_out ),
       .io_VwirePorts_1_13_1_in( ArrayRowModule_1_io_V_wire_out_209 ),
       .io_VwirePorts_1_13_1_en( T577 ),
       .io_VwirePorts_1_13_1_out( VwireModule_io_VwirePorts_1_13_1_out ),
       .io_VwirePorts_1_13_0_in( ArrayRowModule_1_io_V_wire_out_208 ),
       .io_VwirePorts_1_13_0_en( T576 ),
       .io_VwirePorts_1_13_0_out( VwireModule_io_VwirePorts_1_13_0_out ),
       .io_VwirePorts_1_12_15_in( ArrayRowModule_1_io_V_wire_out_207 ),
       .io_VwirePorts_1_12_15_en( T575 ),
       .io_VwirePorts_1_12_15_out( VwireModule_io_VwirePorts_1_12_15_out ),
       .io_VwirePorts_1_12_14_in( ArrayRowModule_1_io_V_wire_out_206 ),
       .io_VwirePorts_1_12_14_en( T574 ),
       .io_VwirePorts_1_12_14_out( VwireModule_io_VwirePorts_1_12_14_out ),
       .io_VwirePorts_1_12_13_in( ArrayRowModule_1_io_V_wire_out_205 ),
       .io_VwirePorts_1_12_13_en( T573 ),
       .io_VwirePorts_1_12_13_out( VwireModule_io_VwirePorts_1_12_13_out ),
       .io_VwirePorts_1_12_12_in( ArrayRowModule_1_io_V_wire_out_204 ),
       .io_VwirePorts_1_12_12_en( T572 ),
       .io_VwirePorts_1_12_12_out( VwireModule_io_VwirePorts_1_12_12_out ),
       .io_VwirePorts_1_12_11_in( ArrayRowModule_1_io_V_wire_out_203 ),
       .io_VwirePorts_1_12_11_en( T571 ),
       .io_VwirePorts_1_12_11_out( VwireModule_io_VwirePorts_1_12_11_out ),
       .io_VwirePorts_1_12_10_in( ArrayRowModule_1_io_V_wire_out_202 ),
       .io_VwirePorts_1_12_10_en( T570 ),
       .io_VwirePorts_1_12_10_out( VwireModule_io_VwirePorts_1_12_10_out ),
       .io_VwirePorts_1_12_9_in( ArrayRowModule_1_io_V_wire_out_201 ),
       .io_VwirePorts_1_12_9_en( T569 ),
       .io_VwirePorts_1_12_9_out( VwireModule_io_VwirePorts_1_12_9_out ),
       .io_VwirePorts_1_12_8_in( ArrayRowModule_1_io_V_wire_out_200 ),
       .io_VwirePorts_1_12_8_en( T568 ),
       .io_VwirePorts_1_12_8_out( VwireModule_io_VwirePorts_1_12_8_out ),
       .io_VwirePorts_1_12_7_in( ArrayRowModule_1_io_V_wire_out_199 ),
       .io_VwirePorts_1_12_7_en( T567 ),
       .io_VwirePorts_1_12_7_out( VwireModule_io_VwirePorts_1_12_7_out ),
       .io_VwirePorts_1_12_6_in( ArrayRowModule_1_io_V_wire_out_198 ),
       .io_VwirePorts_1_12_6_en( T566 ),
       .io_VwirePorts_1_12_6_out( VwireModule_io_VwirePorts_1_12_6_out ),
       .io_VwirePorts_1_12_5_in( ArrayRowModule_1_io_V_wire_out_197 ),
       .io_VwirePorts_1_12_5_en( T565 ),
       .io_VwirePorts_1_12_5_out( VwireModule_io_VwirePorts_1_12_5_out ),
       .io_VwirePorts_1_12_4_in( ArrayRowModule_1_io_V_wire_out_196 ),
       .io_VwirePorts_1_12_4_en( T564 ),
       .io_VwirePorts_1_12_4_out( VwireModule_io_VwirePorts_1_12_4_out ),
       .io_VwirePorts_1_12_3_in( ArrayRowModule_1_io_V_wire_out_195 ),
       .io_VwirePorts_1_12_3_en( T563 ),
       .io_VwirePorts_1_12_3_out( VwireModule_io_VwirePorts_1_12_3_out ),
       .io_VwirePorts_1_12_2_in( ArrayRowModule_1_io_V_wire_out_194 ),
       .io_VwirePorts_1_12_2_en( T562 ),
       .io_VwirePorts_1_12_2_out( VwireModule_io_VwirePorts_1_12_2_out ),
       .io_VwirePorts_1_12_1_in( ArrayRowModule_1_io_V_wire_out_193 ),
       .io_VwirePorts_1_12_1_en( T561 ),
       .io_VwirePorts_1_12_1_out( VwireModule_io_VwirePorts_1_12_1_out ),
       .io_VwirePorts_1_12_0_in( ArrayRowModule_1_io_V_wire_out_192 ),
       .io_VwirePorts_1_12_0_en( T560 ),
       .io_VwirePorts_1_12_0_out( VwireModule_io_VwirePorts_1_12_0_out ),
       .io_VwirePorts_1_11_15_in( ArrayRowModule_1_io_V_wire_out_191 ),
       .io_VwirePorts_1_11_15_en( T559 ),
       .io_VwirePorts_1_11_15_out( VwireModule_io_VwirePorts_1_11_15_out ),
       .io_VwirePorts_1_11_14_in( ArrayRowModule_1_io_V_wire_out_190 ),
       .io_VwirePorts_1_11_14_en( T558 ),
       .io_VwirePorts_1_11_14_out( VwireModule_io_VwirePorts_1_11_14_out ),
       .io_VwirePorts_1_11_13_in( ArrayRowModule_1_io_V_wire_out_189 ),
       .io_VwirePorts_1_11_13_en( T557 ),
       .io_VwirePorts_1_11_13_out( VwireModule_io_VwirePorts_1_11_13_out ),
       .io_VwirePorts_1_11_12_in( ArrayRowModule_1_io_V_wire_out_188 ),
       .io_VwirePorts_1_11_12_en( T556 ),
       .io_VwirePorts_1_11_12_out( VwireModule_io_VwirePorts_1_11_12_out ),
       .io_VwirePorts_1_11_11_in( ArrayRowModule_1_io_V_wire_out_187 ),
       .io_VwirePorts_1_11_11_en( T555 ),
       .io_VwirePorts_1_11_11_out( VwireModule_io_VwirePorts_1_11_11_out ),
       .io_VwirePorts_1_11_10_in( ArrayRowModule_1_io_V_wire_out_186 ),
       .io_VwirePorts_1_11_10_en( T554 ),
       .io_VwirePorts_1_11_10_out( VwireModule_io_VwirePorts_1_11_10_out ),
       .io_VwirePorts_1_11_9_in( ArrayRowModule_1_io_V_wire_out_185 ),
       .io_VwirePorts_1_11_9_en( T553 ),
       .io_VwirePorts_1_11_9_out( VwireModule_io_VwirePorts_1_11_9_out ),
       .io_VwirePorts_1_11_8_in( ArrayRowModule_1_io_V_wire_out_184 ),
       .io_VwirePorts_1_11_8_en( T552 ),
       .io_VwirePorts_1_11_8_out( VwireModule_io_VwirePorts_1_11_8_out ),
       .io_VwirePorts_1_11_7_in( ArrayRowModule_1_io_V_wire_out_183 ),
       .io_VwirePorts_1_11_7_en( T551 ),
       .io_VwirePorts_1_11_7_out( VwireModule_io_VwirePorts_1_11_7_out ),
       .io_VwirePorts_1_11_6_in( ArrayRowModule_1_io_V_wire_out_182 ),
       .io_VwirePorts_1_11_6_en( T550 ),
       .io_VwirePorts_1_11_6_out( VwireModule_io_VwirePorts_1_11_6_out ),
       .io_VwirePorts_1_11_5_in( ArrayRowModule_1_io_V_wire_out_181 ),
       .io_VwirePorts_1_11_5_en( T549 ),
       .io_VwirePorts_1_11_5_out( VwireModule_io_VwirePorts_1_11_5_out ),
       .io_VwirePorts_1_11_4_in( ArrayRowModule_1_io_V_wire_out_180 ),
       .io_VwirePorts_1_11_4_en( T548 ),
       .io_VwirePorts_1_11_4_out( VwireModule_io_VwirePorts_1_11_4_out ),
       .io_VwirePorts_1_11_3_in( ArrayRowModule_1_io_V_wire_out_179 ),
       .io_VwirePorts_1_11_3_en( T547 ),
       .io_VwirePorts_1_11_3_out( VwireModule_io_VwirePorts_1_11_3_out ),
       .io_VwirePorts_1_11_2_in( ArrayRowModule_1_io_V_wire_out_178 ),
       .io_VwirePorts_1_11_2_en( T546 ),
       .io_VwirePorts_1_11_2_out( VwireModule_io_VwirePorts_1_11_2_out ),
       .io_VwirePorts_1_11_1_in( ArrayRowModule_1_io_V_wire_out_177 ),
       .io_VwirePorts_1_11_1_en( T545 ),
       .io_VwirePorts_1_11_1_out( VwireModule_io_VwirePorts_1_11_1_out ),
       .io_VwirePorts_1_11_0_in( ArrayRowModule_1_io_V_wire_out_176 ),
       .io_VwirePorts_1_11_0_en( T544 ),
       .io_VwirePorts_1_11_0_out( VwireModule_io_VwirePorts_1_11_0_out ),
       .io_VwirePorts_1_10_15_in( ArrayRowModule_1_io_V_wire_out_175 ),
       .io_VwirePorts_1_10_15_en( T543 ),
       .io_VwirePorts_1_10_15_out( VwireModule_io_VwirePorts_1_10_15_out ),
       .io_VwirePorts_1_10_14_in( ArrayRowModule_1_io_V_wire_out_174 ),
       .io_VwirePorts_1_10_14_en( T542 ),
       .io_VwirePorts_1_10_14_out( VwireModule_io_VwirePorts_1_10_14_out ),
       .io_VwirePorts_1_10_13_in( ArrayRowModule_1_io_V_wire_out_173 ),
       .io_VwirePorts_1_10_13_en( T541 ),
       .io_VwirePorts_1_10_13_out( VwireModule_io_VwirePorts_1_10_13_out ),
       .io_VwirePorts_1_10_12_in( ArrayRowModule_1_io_V_wire_out_172 ),
       .io_VwirePorts_1_10_12_en( T540 ),
       .io_VwirePorts_1_10_12_out( VwireModule_io_VwirePorts_1_10_12_out ),
       .io_VwirePorts_1_10_11_in( ArrayRowModule_1_io_V_wire_out_171 ),
       .io_VwirePorts_1_10_11_en( T539 ),
       .io_VwirePorts_1_10_11_out( VwireModule_io_VwirePorts_1_10_11_out ),
       .io_VwirePorts_1_10_10_in( ArrayRowModule_1_io_V_wire_out_170 ),
       .io_VwirePorts_1_10_10_en( T538 ),
       .io_VwirePorts_1_10_10_out( VwireModule_io_VwirePorts_1_10_10_out ),
       .io_VwirePorts_1_10_9_in( ArrayRowModule_1_io_V_wire_out_169 ),
       .io_VwirePorts_1_10_9_en( T537 ),
       .io_VwirePorts_1_10_9_out( VwireModule_io_VwirePorts_1_10_9_out ),
       .io_VwirePorts_1_10_8_in( ArrayRowModule_1_io_V_wire_out_168 ),
       .io_VwirePorts_1_10_8_en( T536 ),
       .io_VwirePorts_1_10_8_out( VwireModule_io_VwirePorts_1_10_8_out ),
       .io_VwirePorts_1_10_7_in( ArrayRowModule_1_io_V_wire_out_167 ),
       .io_VwirePorts_1_10_7_en( T535 ),
       .io_VwirePorts_1_10_7_out( VwireModule_io_VwirePorts_1_10_7_out ),
       .io_VwirePorts_1_10_6_in( ArrayRowModule_1_io_V_wire_out_166 ),
       .io_VwirePorts_1_10_6_en( T534 ),
       .io_VwirePorts_1_10_6_out( VwireModule_io_VwirePorts_1_10_6_out ),
       .io_VwirePorts_1_10_5_in( ArrayRowModule_1_io_V_wire_out_165 ),
       .io_VwirePorts_1_10_5_en( T533 ),
       .io_VwirePorts_1_10_5_out( VwireModule_io_VwirePorts_1_10_5_out ),
       .io_VwirePorts_1_10_4_in( ArrayRowModule_1_io_V_wire_out_164 ),
       .io_VwirePorts_1_10_4_en( T532 ),
       .io_VwirePorts_1_10_4_out( VwireModule_io_VwirePorts_1_10_4_out ),
       .io_VwirePorts_1_10_3_in( ArrayRowModule_1_io_V_wire_out_163 ),
       .io_VwirePorts_1_10_3_en( T531 ),
       .io_VwirePorts_1_10_3_out( VwireModule_io_VwirePorts_1_10_3_out ),
       .io_VwirePorts_1_10_2_in( ArrayRowModule_1_io_V_wire_out_162 ),
       .io_VwirePorts_1_10_2_en( T530 ),
       .io_VwirePorts_1_10_2_out( VwireModule_io_VwirePorts_1_10_2_out ),
       .io_VwirePorts_1_10_1_in( ArrayRowModule_1_io_V_wire_out_161 ),
       .io_VwirePorts_1_10_1_en( T529 ),
       .io_VwirePorts_1_10_1_out( VwireModule_io_VwirePorts_1_10_1_out ),
       .io_VwirePorts_1_10_0_in( ArrayRowModule_1_io_V_wire_out_160 ),
       .io_VwirePorts_1_10_0_en( T528 ),
       .io_VwirePorts_1_10_0_out( VwireModule_io_VwirePorts_1_10_0_out ),
       .io_VwirePorts_1_9_15_in( ArrayRowModule_1_io_V_wire_out_159 ),
       .io_VwirePorts_1_9_15_en( T527 ),
       .io_VwirePorts_1_9_15_out( VwireModule_io_VwirePorts_1_9_15_out ),
       .io_VwirePorts_1_9_14_in( ArrayRowModule_1_io_V_wire_out_158 ),
       .io_VwirePorts_1_9_14_en( T526 ),
       .io_VwirePorts_1_9_14_out( VwireModule_io_VwirePorts_1_9_14_out ),
       .io_VwirePorts_1_9_13_in( ArrayRowModule_1_io_V_wire_out_157 ),
       .io_VwirePorts_1_9_13_en( T525 ),
       .io_VwirePorts_1_9_13_out( VwireModule_io_VwirePorts_1_9_13_out ),
       .io_VwirePorts_1_9_12_in( ArrayRowModule_1_io_V_wire_out_156 ),
       .io_VwirePorts_1_9_12_en( T524 ),
       .io_VwirePorts_1_9_12_out( VwireModule_io_VwirePorts_1_9_12_out ),
       .io_VwirePorts_1_9_11_in( ArrayRowModule_1_io_V_wire_out_155 ),
       .io_VwirePorts_1_9_11_en( T523 ),
       .io_VwirePorts_1_9_11_out( VwireModule_io_VwirePorts_1_9_11_out ),
       .io_VwirePorts_1_9_10_in( ArrayRowModule_1_io_V_wire_out_154 ),
       .io_VwirePorts_1_9_10_en( T522 ),
       .io_VwirePorts_1_9_10_out( VwireModule_io_VwirePorts_1_9_10_out ),
       .io_VwirePorts_1_9_9_in( ArrayRowModule_1_io_V_wire_out_153 ),
       .io_VwirePorts_1_9_9_en( T521 ),
       .io_VwirePorts_1_9_9_out( VwireModule_io_VwirePorts_1_9_9_out ),
       .io_VwirePorts_1_9_8_in( ArrayRowModule_1_io_V_wire_out_152 ),
       .io_VwirePorts_1_9_8_en( T520 ),
       .io_VwirePorts_1_9_8_out( VwireModule_io_VwirePorts_1_9_8_out ),
       .io_VwirePorts_1_9_7_in( ArrayRowModule_1_io_V_wire_out_151 ),
       .io_VwirePorts_1_9_7_en( T519 ),
       .io_VwirePorts_1_9_7_out( VwireModule_io_VwirePorts_1_9_7_out ),
       .io_VwirePorts_1_9_6_in( ArrayRowModule_1_io_V_wire_out_150 ),
       .io_VwirePorts_1_9_6_en( T518 ),
       .io_VwirePorts_1_9_6_out( VwireModule_io_VwirePorts_1_9_6_out ),
       .io_VwirePorts_1_9_5_in( ArrayRowModule_1_io_V_wire_out_149 ),
       .io_VwirePorts_1_9_5_en( T517 ),
       .io_VwirePorts_1_9_5_out( VwireModule_io_VwirePorts_1_9_5_out ),
       .io_VwirePorts_1_9_4_in( ArrayRowModule_1_io_V_wire_out_148 ),
       .io_VwirePorts_1_9_4_en( T516 ),
       .io_VwirePorts_1_9_4_out( VwireModule_io_VwirePorts_1_9_4_out ),
       .io_VwirePorts_1_9_3_in( ArrayRowModule_1_io_V_wire_out_147 ),
       .io_VwirePorts_1_9_3_en( T515 ),
       .io_VwirePorts_1_9_3_out( VwireModule_io_VwirePorts_1_9_3_out ),
       .io_VwirePorts_1_9_2_in( ArrayRowModule_1_io_V_wire_out_146 ),
       .io_VwirePorts_1_9_2_en( T514 ),
       .io_VwirePorts_1_9_2_out( VwireModule_io_VwirePorts_1_9_2_out ),
       .io_VwirePorts_1_9_1_in( ArrayRowModule_1_io_V_wire_out_145 ),
       .io_VwirePorts_1_9_1_en( T513 ),
       .io_VwirePorts_1_9_1_out( VwireModule_io_VwirePorts_1_9_1_out ),
       .io_VwirePorts_1_9_0_in( ArrayRowModule_1_io_V_wire_out_144 ),
       .io_VwirePorts_1_9_0_en( T512 ),
       .io_VwirePorts_1_9_0_out( VwireModule_io_VwirePorts_1_9_0_out ),
       .io_VwirePorts_1_8_15_in( ArrayRowModule_1_io_V_wire_out_143 ),
       .io_VwirePorts_1_8_15_en( T511 ),
       .io_VwirePorts_1_8_15_out( VwireModule_io_VwirePorts_1_8_15_out ),
       .io_VwirePorts_1_8_14_in( ArrayRowModule_1_io_V_wire_out_142 ),
       .io_VwirePorts_1_8_14_en( T510 ),
       .io_VwirePorts_1_8_14_out( VwireModule_io_VwirePorts_1_8_14_out ),
       .io_VwirePorts_1_8_13_in( ArrayRowModule_1_io_V_wire_out_141 ),
       .io_VwirePorts_1_8_13_en( T509 ),
       .io_VwirePorts_1_8_13_out( VwireModule_io_VwirePorts_1_8_13_out ),
       .io_VwirePorts_1_8_12_in( ArrayRowModule_1_io_V_wire_out_140 ),
       .io_VwirePorts_1_8_12_en( T508 ),
       .io_VwirePorts_1_8_12_out( VwireModule_io_VwirePorts_1_8_12_out ),
       .io_VwirePorts_1_8_11_in( ArrayRowModule_1_io_V_wire_out_139 ),
       .io_VwirePorts_1_8_11_en( T507 ),
       .io_VwirePorts_1_8_11_out( VwireModule_io_VwirePorts_1_8_11_out ),
       .io_VwirePorts_1_8_10_in( ArrayRowModule_1_io_V_wire_out_138 ),
       .io_VwirePorts_1_8_10_en( T506 ),
       .io_VwirePorts_1_8_10_out( VwireModule_io_VwirePorts_1_8_10_out ),
       .io_VwirePorts_1_8_9_in( ArrayRowModule_1_io_V_wire_out_137 ),
       .io_VwirePorts_1_8_9_en( T505 ),
       .io_VwirePorts_1_8_9_out( VwireModule_io_VwirePorts_1_8_9_out ),
       .io_VwirePorts_1_8_8_in( ArrayRowModule_1_io_V_wire_out_136 ),
       .io_VwirePorts_1_8_8_en( T504 ),
       .io_VwirePorts_1_8_8_out( VwireModule_io_VwirePorts_1_8_8_out ),
       .io_VwirePorts_1_8_7_in( ArrayRowModule_1_io_V_wire_out_135 ),
       .io_VwirePorts_1_8_7_en( T503 ),
       .io_VwirePorts_1_8_7_out( VwireModule_io_VwirePorts_1_8_7_out ),
       .io_VwirePorts_1_8_6_in( ArrayRowModule_1_io_V_wire_out_134 ),
       .io_VwirePorts_1_8_6_en( T502 ),
       .io_VwirePorts_1_8_6_out( VwireModule_io_VwirePorts_1_8_6_out ),
       .io_VwirePorts_1_8_5_in( ArrayRowModule_1_io_V_wire_out_133 ),
       .io_VwirePorts_1_8_5_en( T501 ),
       .io_VwirePorts_1_8_5_out( VwireModule_io_VwirePorts_1_8_5_out ),
       .io_VwirePorts_1_8_4_in( ArrayRowModule_1_io_V_wire_out_132 ),
       .io_VwirePorts_1_8_4_en( T500 ),
       .io_VwirePorts_1_8_4_out( VwireModule_io_VwirePorts_1_8_4_out ),
       .io_VwirePorts_1_8_3_in( ArrayRowModule_1_io_V_wire_out_131 ),
       .io_VwirePorts_1_8_3_en( T499 ),
       .io_VwirePorts_1_8_3_out( VwireModule_io_VwirePorts_1_8_3_out ),
       .io_VwirePorts_1_8_2_in( ArrayRowModule_1_io_V_wire_out_130 ),
       .io_VwirePorts_1_8_2_en( T498 ),
       .io_VwirePorts_1_8_2_out( VwireModule_io_VwirePorts_1_8_2_out ),
       .io_VwirePorts_1_8_1_in( ArrayRowModule_1_io_V_wire_out_129 ),
       .io_VwirePorts_1_8_1_en( T497 ),
       .io_VwirePorts_1_8_1_out( VwireModule_io_VwirePorts_1_8_1_out ),
       .io_VwirePorts_1_8_0_in( ArrayRowModule_1_io_V_wire_out_128 ),
       .io_VwirePorts_1_8_0_en( T496 ),
       .io_VwirePorts_1_8_0_out( VwireModule_io_VwirePorts_1_8_0_out ),
       .io_VwirePorts_1_7_15_in( ArrayRowModule_1_io_V_wire_out_127 ),
       .io_VwirePorts_1_7_15_en( T495 ),
       .io_VwirePorts_1_7_15_out( VwireModule_io_VwirePorts_1_7_15_out ),
       .io_VwirePorts_1_7_14_in( ArrayRowModule_1_io_V_wire_out_126 ),
       .io_VwirePorts_1_7_14_en( T494 ),
       .io_VwirePorts_1_7_14_out( VwireModule_io_VwirePorts_1_7_14_out ),
       .io_VwirePorts_1_7_13_in( ArrayRowModule_1_io_V_wire_out_125 ),
       .io_VwirePorts_1_7_13_en( T493 ),
       .io_VwirePorts_1_7_13_out( VwireModule_io_VwirePorts_1_7_13_out ),
       .io_VwirePorts_1_7_12_in( ArrayRowModule_1_io_V_wire_out_124 ),
       .io_VwirePorts_1_7_12_en( T492 ),
       .io_VwirePorts_1_7_12_out( VwireModule_io_VwirePorts_1_7_12_out ),
       .io_VwirePorts_1_7_11_in( ArrayRowModule_1_io_V_wire_out_123 ),
       .io_VwirePorts_1_7_11_en( T491 ),
       .io_VwirePorts_1_7_11_out( VwireModule_io_VwirePorts_1_7_11_out ),
       .io_VwirePorts_1_7_10_in( ArrayRowModule_1_io_V_wire_out_122 ),
       .io_VwirePorts_1_7_10_en( T490 ),
       .io_VwirePorts_1_7_10_out( VwireModule_io_VwirePorts_1_7_10_out ),
       .io_VwirePorts_1_7_9_in( ArrayRowModule_1_io_V_wire_out_121 ),
       .io_VwirePorts_1_7_9_en( T489 ),
       .io_VwirePorts_1_7_9_out( VwireModule_io_VwirePorts_1_7_9_out ),
       .io_VwirePorts_1_7_8_in( ArrayRowModule_1_io_V_wire_out_120 ),
       .io_VwirePorts_1_7_8_en( T488 ),
       .io_VwirePorts_1_7_8_out( VwireModule_io_VwirePorts_1_7_8_out ),
       .io_VwirePorts_1_7_7_in( ArrayRowModule_1_io_V_wire_out_119 ),
       .io_VwirePorts_1_7_7_en( T487 ),
       .io_VwirePorts_1_7_7_out( VwireModule_io_VwirePorts_1_7_7_out ),
       .io_VwirePorts_1_7_6_in( ArrayRowModule_1_io_V_wire_out_118 ),
       .io_VwirePorts_1_7_6_en( T486 ),
       .io_VwirePorts_1_7_6_out( VwireModule_io_VwirePorts_1_7_6_out ),
       .io_VwirePorts_1_7_5_in( ArrayRowModule_1_io_V_wire_out_117 ),
       .io_VwirePorts_1_7_5_en( T485 ),
       .io_VwirePorts_1_7_5_out( VwireModule_io_VwirePorts_1_7_5_out ),
       .io_VwirePorts_1_7_4_in( ArrayRowModule_1_io_V_wire_out_116 ),
       .io_VwirePorts_1_7_4_en( T484 ),
       .io_VwirePorts_1_7_4_out( VwireModule_io_VwirePorts_1_7_4_out ),
       .io_VwirePorts_1_7_3_in( ArrayRowModule_1_io_V_wire_out_115 ),
       .io_VwirePorts_1_7_3_en( T483 ),
       .io_VwirePorts_1_7_3_out( VwireModule_io_VwirePorts_1_7_3_out ),
       .io_VwirePorts_1_7_2_in( ArrayRowModule_1_io_V_wire_out_114 ),
       .io_VwirePorts_1_7_2_en( T482 ),
       .io_VwirePorts_1_7_2_out( VwireModule_io_VwirePorts_1_7_2_out ),
       .io_VwirePorts_1_7_1_in( ArrayRowModule_1_io_V_wire_out_113 ),
       .io_VwirePorts_1_7_1_en( T481 ),
       .io_VwirePorts_1_7_1_out( VwireModule_io_VwirePorts_1_7_1_out ),
       .io_VwirePorts_1_7_0_in( ArrayRowModule_1_io_V_wire_out_112 ),
       .io_VwirePorts_1_7_0_en( T480 ),
       .io_VwirePorts_1_7_0_out( VwireModule_io_VwirePorts_1_7_0_out ),
       .io_VwirePorts_1_6_15_in( ArrayRowModule_1_io_V_wire_out_111 ),
       .io_VwirePorts_1_6_15_en( T479 ),
       .io_VwirePorts_1_6_15_out( VwireModule_io_VwirePorts_1_6_15_out ),
       .io_VwirePorts_1_6_14_in( ArrayRowModule_1_io_V_wire_out_110 ),
       .io_VwirePorts_1_6_14_en( T478 ),
       .io_VwirePorts_1_6_14_out( VwireModule_io_VwirePorts_1_6_14_out ),
       .io_VwirePorts_1_6_13_in( ArrayRowModule_1_io_V_wire_out_109 ),
       .io_VwirePorts_1_6_13_en( T477 ),
       .io_VwirePorts_1_6_13_out( VwireModule_io_VwirePorts_1_6_13_out ),
       .io_VwirePorts_1_6_12_in( ArrayRowModule_1_io_V_wire_out_108 ),
       .io_VwirePorts_1_6_12_en( T476 ),
       .io_VwirePorts_1_6_12_out( VwireModule_io_VwirePorts_1_6_12_out ),
       .io_VwirePorts_1_6_11_in( ArrayRowModule_1_io_V_wire_out_107 ),
       .io_VwirePorts_1_6_11_en( T475 ),
       .io_VwirePorts_1_6_11_out( VwireModule_io_VwirePorts_1_6_11_out ),
       .io_VwirePorts_1_6_10_in( ArrayRowModule_1_io_V_wire_out_106 ),
       .io_VwirePorts_1_6_10_en( T474 ),
       .io_VwirePorts_1_6_10_out( VwireModule_io_VwirePorts_1_6_10_out ),
       .io_VwirePorts_1_6_9_in( ArrayRowModule_1_io_V_wire_out_105 ),
       .io_VwirePorts_1_6_9_en( T473 ),
       .io_VwirePorts_1_6_9_out( VwireModule_io_VwirePorts_1_6_9_out ),
       .io_VwirePorts_1_6_8_in( ArrayRowModule_1_io_V_wire_out_104 ),
       .io_VwirePorts_1_6_8_en( T472 ),
       .io_VwirePorts_1_6_8_out( VwireModule_io_VwirePorts_1_6_8_out ),
       .io_VwirePorts_1_6_7_in( ArrayRowModule_1_io_V_wire_out_103 ),
       .io_VwirePorts_1_6_7_en( T471 ),
       .io_VwirePorts_1_6_7_out( VwireModule_io_VwirePorts_1_6_7_out ),
       .io_VwirePorts_1_6_6_in( ArrayRowModule_1_io_V_wire_out_102 ),
       .io_VwirePorts_1_6_6_en( T470 ),
       .io_VwirePorts_1_6_6_out( VwireModule_io_VwirePorts_1_6_6_out ),
       .io_VwirePorts_1_6_5_in( ArrayRowModule_1_io_V_wire_out_101 ),
       .io_VwirePorts_1_6_5_en( T469 ),
       .io_VwirePorts_1_6_5_out( VwireModule_io_VwirePorts_1_6_5_out ),
       .io_VwirePorts_1_6_4_in( ArrayRowModule_1_io_V_wire_out_100 ),
       .io_VwirePorts_1_6_4_en( T468 ),
       .io_VwirePorts_1_6_4_out( VwireModule_io_VwirePorts_1_6_4_out ),
       .io_VwirePorts_1_6_3_in( ArrayRowModule_1_io_V_wire_out_99 ),
       .io_VwirePorts_1_6_3_en( T467 ),
       .io_VwirePorts_1_6_3_out( VwireModule_io_VwirePorts_1_6_3_out ),
       .io_VwirePorts_1_6_2_in( ArrayRowModule_1_io_V_wire_out_98 ),
       .io_VwirePorts_1_6_2_en( T466 ),
       .io_VwirePorts_1_6_2_out( VwireModule_io_VwirePorts_1_6_2_out ),
       .io_VwirePorts_1_6_1_in( ArrayRowModule_1_io_V_wire_out_97 ),
       .io_VwirePorts_1_6_1_en( T465 ),
       .io_VwirePorts_1_6_1_out( VwireModule_io_VwirePorts_1_6_1_out ),
       .io_VwirePorts_1_6_0_in( ArrayRowModule_1_io_V_wire_out_96 ),
       .io_VwirePorts_1_6_0_en( T464 ),
       .io_VwirePorts_1_6_0_out( VwireModule_io_VwirePorts_1_6_0_out ),
       .io_VwirePorts_1_5_15_in( ArrayRowModule_1_io_V_wire_out_95 ),
       .io_VwirePorts_1_5_15_en( T463 ),
       .io_VwirePorts_1_5_15_out( VwireModule_io_VwirePorts_1_5_15_out ),
       .io_VwirePorts_1_5_14_in( ArrayRowModule_1_io_V_wire_out_94 ),
       .io_VwirePorts_1_5_14_en( T462 ),
       .io_VwirePorts_1_5_14_out( VwireModule_io_VwirePorts_1_5_14_out ),
       .io_VwirePorts_1_5_13_in( ArrayRowModule_1_io_V_wire_out_93 ),
       .io_VwirePorts_1_5_13_en( T461 ),
       .io_VwirePorts_1_5_13_out( VwireModule_io_VwirePorts_1_5_13_out ),
       .io_VwirePorts_1_5_12_in( ArrayRowModule_1_io_V_wire_out_92 ),
       .io_VwirePorts_1_5_12_en( T460 ),
       .io_VwirePorts_1_5_12_out( VwireModule_io_VwirePorts_1_5_12_out ),
       .io_VwirePorts_1_5_11_in( ArrayRowModule_1_io_V_wire_out_91 ),
       .io_VwirePorts_1_5_11_en( T459 ),
       .io_VwirePorts_1_5_11_out( VwireModule_io_VwirePorts_1_5_11_out ),
       .io_VwirePorts_1_5_10_in( ArrayRowModule_1_io_V_wire_out_90 ),
       .io_VwirePorts_1_5_10_en( T458 ),
       .io_VwirePorts_1_5_10_out( VwireModule_io_VwirePorts_1_5_10_out ),
       .io_VwirePorts_1_5_9_in( ArrayRowModule_1_io_V_wire_out_89 ),
       .io_VwirePorts_1_5_9_en( T457 ),
       .io_VwirePorts_1_5_9_out( VwireModule_io_VwirePorts_1_5_9_out ),
       .io_VwirePorts_1_5_8_in( ArrayRowModule_1_io_V_wire_out_88 ),
       .io_VwirePorts_1_5_8_en( T456 ),
       .io_VwirePorts_1_5_8_out( VwireModule_io_VwirePorts_1_5_8_out ),
       .io_VwirePorts_1_5_7_in( ArrayRowModule_1_io_V_wire_out_87 ),
       .io_VwirePorts_1_5_7_en( T455 ),
       .io_VwirePorts_1_5_7_out( VwireModule_io_VwirePorts_1_5_7_out ),
       .io_VwirePorts_1_5_6_in( ArrayRowModule_1_io_V_wire_out_86 ),
       .io_VwirePorts_1_5_6_en( T454 ),
       .io_VwirePorts_1_5_6_out( VwireModule_io_VwirePorts_1_5_6_out ),
       .io_VwirePorts_1_5_5_in( ArrayRowModule_1_io_V_wire_out_85 ),
       .io_VwirePorts_1_5_5_en( T453 ),
       .io_VwirePorts_1_5_5_out( VwireModule_io_VwirePorts_1_5_5_out ),
       .io_VwirePorts_1_5_4_in( ArrayRowModule_1_io_V_wire_out_84 ),
       .io_VwirePorts_1_5_4_en( T452 ),
       .io_VwirePorts_1_5_4_out( VwireModule_io_VwirePorts_1_5_4_out ),
       .io_VwirePorts_1_5_3_in( ArrayRowModule_1_io_V_wire_out_83 ),
       .io_VwirePorts_1_5_3_en( T451 ),
       .io_VwirePorts_1_5_3_out( VwireModule_io_VwirePorts_1_5_3_out ),
       .io_VwirePorts_1_5_2_in( ArrayRowModule_1_io_V_wire_out_82 ),
       .io_VwirePorts_1_5_2_en( T450 ),
       .io_VwirePorts_1_5_2_out( VwireModule_io_VwirePorts_1_5_2_out ),
       .io_VwirePorts_1_5_1_in( ArrayRowModule_1_io_V_wire_out_81 ),
       .io_VwirePorts_1_5_1_en( T449 ),
       .io_VwirePorts_1_5_1_out( VwireModule_io_VwirePorts_1_5_1_out ),
       .io_VwirePorts_1_5_0_in( ArrayRowModule_1_io_V_wire_out_80 ),
       .io_VwirePorts_1_5_0_en( T448 ),
       .io_VwirePorts_1_5_0_out( VwireModule_io_VwirePorts_1_5_0_out ),
       .io_VwirePorts_1_4_15_in( ArrayRowModule_1_io_V_wire_out_79 ),
       .io_VwirePorts_1_4_15_en( T447 ),
       .io_VwirePorts_1_4_15_out( VwireModule_io_VwirePorts_1_4_15_out ),
       .io_VwirePorts_1_4_14_in( ArrayRowModule_1_io_V_wire_out_78 ),
       .io_VwirePorts_1_4_14_en( T446 ),
       .io_VwirePorts_1_4_14_out( VwireModule_io_VwirePorts_1_4_14_out ),
       .io_VwirePorts_1_4_13_in( ArrayRowModule_1_io_V_wire_out_77 ),
       .io_VwirePorts_1_4_13_en( T445 ),
       .io_VwirePorts_1_4_13_out( VwireModule_io_VwirePorts_1_4_13_out ),
       .io_VwirePorts_1_4_12_in( ArrayRowModule_1_io_V_wire_out_76 ),
       .io_VwirePorts_1_4_12_en( T444 ),
       .io_VwirePorts_1_4_12_out( VwireModule_io_VwirePorts_1_4_12_out ),
       .io_VwirePorts_1_4_11_in( ArrayRowModule_1_io_V_wire_out_75 ),
       .io_VwirePorts_1_4_11_en( T443 ),
       .io_VwirePorts_1_4_11_out( VwireModule_io_VwirePorts_1_4_11_out ),
       .io_VwirePorts_1_4_10_in( ArrayRowModule_1_io_V_wire_out_74 ),
       .io_VwirePorts_1_4_10_en( T442 ),
       .io_VwirePorts_1_4_10_out( VwireModule_io_VwirePorts_1_4_10_out ),
       .io_VwirePorts_1_4_9_in( ArrayRowModule_1_io_V_wire_out_73 ),
       .io_VwirePorts_1_4_9_en( T441 ),
       .io_VwirePorts_1_4_9_out( VwireModule_io_VwirePorts_1_4_9_out ),
       .io_VwirePorts_1_4_8_in( ArrayRowModule_1_io_V_wire_out_72 ),
       .io_VwirePorts_1_4_8_en( T440 ),
       .io_VwirePorts_1_4_8_out( VwireModule_io_VwirePorts_1_4_8_out ),
       .io_VwirePorts_1_4_7_in( ArrayRowModule_1_io_V_wire_out_71 ),
       .io_VwirePorts_1_4_7_en( T439 ),
       .io_VwirePorts_1_4_7_out( VwireModule_io_VwirePorts_1_4_7_out ),
       .io_VwirePorts_1_4_6_in( ArrayRowModule_1_io_V_wire_out_70 ),
       .io_VwirePorts_1_4_6_en( T438 ),
       .io_VwirePorts_1_4_6_out( VwireModule_io_VwirePorts_1_4_6_out ),
       .io_VwirePorts_1_4_5_in( ArrayRowModule_1_io_V_wire_out_69 ),
       .io_VwirePorts_1_4_5_en( T437 ),
       .io_VwirePorts_1_4_5_out( VwireModule_io_VwirePorts_1_4_5_out ),
       .io_VwirePorts_1_4_4_in( ArrayRowModule_1_io_V_wire_out_68 ),
       .io_VwirePorts_1_4_4_en( T436 ),
       .io_VwirePorts_1_4_4_out( VwireModule_io_VwirePorts_1_4_4_out ),
       .io_VwirePorts_1_4_3_in( ArrayRowModule_1_io_V_wire_out_67 ),
       .io_VwirePorts_1_4_3_en( T435 ),
       .io_VwirePorts_1_4_3_out( VwireModule_io_VwirePorts_1_4_3_out ),
       .io_VwirePorts_1_4_2_in( ArrayRowModule_1_io_V_wire_out_66 ),
       .io_VwirePorts_1_4_2_en( T434 ),
       .io_VwirePorts_1_4_2_out( VwireModule_io_VwirePorts_1_4_2_out ),
       .io_VwirePorts_1_4_1_in( ArrayRowModule_1_io_V_wire_out_65 ),
       .io_VwirePorts_1_4_1_en( T433 ),
       .io_VwirePorts_1_4_1_out( VwireModule_io_VwirePorts_1_4_1_out ),
       .io_VwirePorts_1_4_0_in( ArrayRowModule_1_io_V_wire_out_64 ),
       .io_VwirePorts_1_4_0_en( T432 ),
       .io_VwirePorts_1_4_0_out( VwireModule_io_VwirePorts_1_4_0_out ),
       .io_VwirePorts_1_3_15_in( ArrayRowModule_1_io_V_wire_out_63 ),
       .io_VwirePorts_1_3_15_en( T431 ),
       .io_VwirePorts_1_3_15_out( VwireModule_io_VwirePorts_1_3_15_out ),
       .io_VwirePorts_1_3_14_in( ArrayRowModule_1_io_V_wire_out_62 ),
       .io_VwirePorts_1_3_14_en( T430 ),
       .io_VwirePorts_1_3_14_out( VwireModule_io_VwirePorts_1_3_14_out ),
       .io_VwirePorts_1_3_13_in( ArrayRowModule_1_io_V_wire_out_61 ),
       .io_VwirePorts_1_3_13_en( T429 ),
       .io_VwirePorts_1_3_13_out( VwireModule_io_VwirePorts_1_3_13_out ),
       .io_VwirePorts_1_3_12_in( ArrayRowModule_1_io_V_wire_out_60 ),
       .io_VwirePorts_1_3_12_en( T428 ),
       .io_VwirePorts_1_3_12_out( VwireModule_io_VwirePorts_1_3_12_out ),
       .io_VwirePorts_1_3_11_in( ArrayRowModule_1_io_V_wire_out_59 ),
       .io_VwirePorts_1_3_11_en( T427 ),
       .io_VwirePorts_1_3_11_out( VwireModule_io_VwirePorts_1_3_11_out ),
       .io_VwirePorts_1_3_10_in( ArrayRowModule_1_io_V_wire_out_58 ),
       .io_VwirePorts_1_3_10_en( T426 ),
       .io_VwirePorts_1_3_10_out( VwireModule_io_VwirePorts_1_3_10_out ),
       .io_VwirePorts_1_3_9_in( ArrayRowModule_1_io_V_wire_out_57 ),
       .io_VwirePorts_1_3_9_en( T425 ),
       .io_VwirePorts_1_3_9_out( VwireModule_io_VwirePorts_1_3_9_out ),
       .io_VwirePorts_1_3_8_in( ArrayRowModule_1_io_V_wire_out_56 ),
       .io_VwirePorts_1_3_8_en( T424 ),
       .io_VwirePorts_1_3_8_out( VwireModule_io_VwirePorts_1_3_8_out ),
       .io_VwirePorts_1_3_7_in( ArrayRowModule_1_io_V_wire_out_55 ),
       .io_VwirePorts_1_3_7_en( T423 ),
       .io_VwirePorts_1_3_7_out( VwireModule_io_VwirePorts_1_3_7_out ),
       .io_VwirePorts_1_3_6_in( ArrayRowModule_1_io_V_wire_out_54 ),
       .io_VwirePorts_1_3_6_en( T422 ),
       .io_VwirePorts_1_3_6_out( VwireModule_io_VwirePorts_1_3_6_out ),
       .io_VwirePorts_1_3_5_in( ArrayRowModule_1_io_V_wire_out_53 ),
       .io_VwirePorts_1_3_5_en( T421 ),
       .io_VwirePorts_1_3_5_out( VwireModule_io_VwirePorts_1_3_5_out ),
       .io_VwirePorts_1_3_4_in( ArrayRowModule_1_io_V_wire_out_52 ),
       .io_VwirePorts_1_3_4_en( T420 ),
       .io_VwirePorts_1_3_4_out( VwireModule_io_VwirePorts_1_3_4_out ),
       .io_VwirePorts_1_3_3_in( ArrayRowModule_1_io_V_wire_out_51 ),
       .io_VwirePorts_1_3_3_en( T419 ),
       .io_VwirePorts_1_3_3_out( VwireModule_io_VwirePorts_1_3_3_out ),
       .io_VwirePorts_1_3_2_in( ArrayRowModule_1_io_V_wire_out_50 ),
       .io_VwirePorts_1_3_2_en( T418 ),
       .io_VwirePorts_1_3_2_out( VwireModule_io_VwirePorts_1_3_2_out ),
       .io_VwirePorts_1_3_1_in( ArrayRowModule_1_io_V_wire_out_49 ),
       .io_VwirePorts_1_3_1_en( T417 ),
       .io_VwirePorts_1_3_1_out( VwireModule_io_VwirePorts_1_3_1_out ),
       .io_VwirePorts_1_3_0_in( ArrayRowModule_1_io_V_wire_out_48 ),
       .io_VwirePorts_1_3_0_en( T416 ),
       .io_VwirePorts_1_3_0_out( VwireModule_io_VwirePorts_1_3_0_out ),
       .io_VwirePorts_1_2_15_in( ArrayRowModule_1_io_V_wire_out_47 ),
       .io_VwirePorts_1_2_15_en( T415 ),
       .io_VwirePorts_1_2_15_out( VwireModule_io_VwirePorts_1_2_15_out ),
       .io_VwirePorts_1_2_14_in( ArrayRowModule_1_io_V_wire_out_46 ),
       .io_VwirePorts_1_2_14_en( T414 ),
       .io_VwirePorts_1_2_14_out( VwireModule_io_VwirePorts_1_2_14_out ),
       .io_VwirePorts_1_2_13_in( ArrayRowModule_1_io_V_wire_out_45 ),
       .io_VwirePorts_1_2_13_en( T413 ),
       .io_VwirePorts_1_2_13_out( VwireModule_io_VwirePorts_1_2_13_out ),
       .io_VwirePorts_1_2_12_in( ArrayRowModule_1_io_V_wire_out_44 ),
       .io_VwirePorts_1_2_12_en( T412 ),
       .io_VwirePorts_1_2_12_out( VwireModule_io_VwirePorts_1_2_12_out ),
       .io_VwirePorts_1_2_11_in( ArrayRowModule_1_io_V_wire_out_43 ),
       .io_VwirePorts_1_2_11_en( T411 ),
       .io_VwirePorts_1_2_11_out( VwireModule_io_VwirePorts_1_2_11_out ),
       .io_VwirePorts_1_2_10_in( ArrayRowModule_1_io_V_wire_out_42 ),
       .io_VwirePorts_1_2_10_en( T410 ),
       .io_VwirePorts_1_2_10_out( VwireModule_io_VwirePorts_1_2_10_out ),
       .io_VwirePorts_1_2_9_in( ArrayRowModule_1_io_V_wire_out_41 ),
       .io_VwirePorts_1_2_9_en( T409 ),
       .io_VwirePorts_1_2_9_out( VwireModule_io_VwirePorts_1_2_9_out ),
       .io_VwirePorts_1_2_8_in( ArrayRowModule_1_io_V_wire_out_40 ),
       .io_VwirePorts_1_2_8_en( T408 ),
       .io_VwirePorts_1_2_8_out( VwireModule_io_VwirePorts_1_2_8_out ),
       .io_VwirePorts_1_2_7_in( ArrayRowModule_1_io_V_wire_out_39 ),
       .io_VwirePorts_1_2_7_en( T407 ),
       .io_VwirePorts_1_2_7_out( VwireModule_io_VwirePorts_1_2_7_out ),
       .io_VwirePorts_1_2_6_in( ArrayRowModule_1_io_V_wire_out_38 ),
       .io_VwirePorts_1_2_6_en( T406 ),
       .io_VwirePorts_1_2_6_out( VwireModule_io_VwirePorts_1_2_6_out ),
       .io_VwirePorts_1_2_5_in( ArrayRowModule_1_io_V_wire_out_37 ),
       .io_VwirePorts_1_2_5_en( T405 ),
       .io_VwirePorts_1_2_5_out( VwireModule_io_VwirePorts_1_2_5_out ),
       .io_VwirePorts_1_2_4_in( ArrayRowModule_1_io_V_wire_out_36 ),
       .io_VwirePorts_1_2_4_en( T404 ),
       .io_VwirePorts_1_2_4_out( VwireModule_io_VwirePorts_1_2_4_out ),
       .io_VwirePorts_1_2_3_in( ArrayRowModule_1_io_V_wire_out_35 ),
       .io_VwirePorts_1_2_3_en( T403 ),
       .io_VwirePorts_1_2_3_out( VwireModule_io_VwirePorts_1_2_3_out ),
       .io_VwirePorts_1_2_2_in( ArrayRowModule_1_io_V_wire_out_34 ),
       .io_VwirePorts_1_2_2_en( T402 ),
       .io_VwirePorts_1_2_2_out( VwireModule_io_VwirePorts_1_2_2_out ),
       .io_VwirePorts_1_2_1_in( ArrayRowModule_1_io_V_wire_out_33 ),
       .io_VwirePorts_1_2_1_en( T401 ),
       .io_VwirePorts_1_2_1_out( VwireModule_io_VwirePorts_1_2_1_out ),
       .io_VwirePorts_1_2_0_in( ArrayRowModule_1_io_V_wire_out_32 ),
       .io_VwirePorts_1_2_0_en( T400 ),
       .io_VwirePorts_1_2_0_out( VwireModule_io_VwirePorts_1_2_0_out ),
       .io_VwirePorts_1_1_15_in( ArrayRowModule_1_io_V_wire_out_31 ),
       .io_VwirePorts_1_1_15_en( T399 ),
       .io_VwirePorts_1_1_15_out( VwireModule_io_VwirePorts_1_1_15_out ),
       .io_VwirePorts_1_1_14_in( ArrayRowModule_1_io_V_wire_out_30 ),
       .io_VwirePorts_1_1_14_en( T398 ),
       .io_VwirePorts_1_1_14_out( VwireModule_io_VwirePorts_1_1_14_out ),
       .io_VwirePorts_1_1_13_in( ArrayRowModule_1_io_V_wire_out_29 ),
       .io_VwirePorts_1_1_13_en( T397 ),
       .io_VwirePorts_1_1_13_out( VwireModule_io_VwirePorts_1_1_13_out ),
       .io_VwirePorts_1_1_12_in( ArrayRowModule_1_io_V_wire_out_28 ),
       .io_VwirePorts_1_1_12_en( T396 ),
       .io_VwirePorts_1_1_12_out( VwireModule_io_VwirePorts_1_1_12_out ),
       .io_VwirePorts_1_1_11_in( ArrayRowModule_1_io_V_wire_out_27 ),
       .io_VwirePorts_1_1_11_en( T395 ),
       .io_VwirePorts_1_1_11_out( VwireModule_io_VwirePorts_1_1_11_out ),
       .io_VwirePorts_1_1_10_in( ArrayRowModule_1_io_V_wire_out_26 ),
       .io_VwirePorts_1_1_10_en( T394 ),
       .io_VwirePorts_1_1_10_out( VwireModule_io_VwirePorts_1_1_10_out ),
       .io_VwirePorts_1_1_9_in( ArrayRowModule_1_io_V_wire_out_25 ),
       .io_VwirePorts_1_1_9_en( T393 ),
       .io_VwirePorts_1_1_9_out( VwireModule_io_VwirePorts_1_1_9_out ),
       .io_VwirePorts_1_1_8_in( ArrayRowModule_1_io_V_wire_out_24 ),
       .io_VwirePorts_1_1_8_en( T392 ),
       .io_VwirePorts_1_1_8_out( VwireModule_io_VwirePorts_1_1_8_out ),
       .io_VwirePorts_1_1_7_in( ArrayRowModule_1_io_V_wire_out_23 ),
       .io_VwirePorts_1_1_7_en( T391 ),
       .io_VwirePorts_1_1_7_out( VwireModule_io_VwirePorts_1_1_7_out ),
       .io_VwirePorts_1_1_6_in( ArrayRowModule_1_io_V_wire_out_22 ),
       .io_VwirePorts_1_1_6_en( T390 ),
       .io_VwirePorts_1_1_6_out( VwireModule_io_VwirePorts_1_1_6_out ),
       .io_VwirePorts_1_1_5_in( ArrayRowModule_1_io_V_wire_out_21 ),
       .io_VwirePorts_1_1_5_en( T389 ),
       .io_VwirePorts_1_1_5_out( VwireModule_io_VwirePorts_1_1_5_out ),
       .io_VwirePorts_1_1_4_in( ArrayRowModule_1_io_V_wire_out_20 ),
       .io_VwirePorts_1_1_4_en( T388 ),
       .io_VwirePorts_1_1_4_out( VwireModule_io_VwirePorts_1_1_4_out ),
       .io_VwirePorts_1_1_3_in( ArrayRowModule_1_io_V_wire_out_19 ),
       .io_VwirePorts_1_1_3_en( T387 ),
       .io_VwirePorts_1_1_3_out( VwireModule_io_VwirePorts_1_1_3_out ),
       .io_VwirePorts_1_1_2_in( ArrayRowModule_1_io_V_wire_out_18 ),
       .io_VwirePorts_1_1_2_en( T386 ),
       .io_VwirePorts_1_1_2_out( VwireModule_io_VwirePorts_1_1_2_out ),
       .io_VwirePorts_1_1_1_in( ArrayRowModule_1_io_V_wire_out_17 ),
       .io_VwirePorts_1_1_1_en( T385 ),
       .io_VwirePorts_1_1_1_out( VwireModule_io_VwirePorts_1_1_1_out ),
       .io_VwirePorts_1_1_0_in( ArrayRowModule_1_io_V_wire_out_16 ),
       .io_VwirePorts_1_1_0_en( T384 ),
       .io_VwirePorts_1_1_0_out( VwireModule_io_VwirePorts_1_1_0_out ),
       .io_VwirePorts_1_0_15_in( ArrayRowModule_1_io_V_wire_out_15 ),
       .io_VwirePorts_1_0_15_en( T383 ),
       .io_VwirePorts_1_0_15_out( VwireModule_io_VwirePorts_1_0_15_out ),
       .io_VwirePorts_1_0_14_in( ArrayRowModule_1_io_V_wire_out_14 ),
       .io_VwirePorts_1_0_14_en( T382 ),
       .io_VwirePorts_1_0_14_out( VwireModule_io_VwirePorts_1_0_14_out ),
       .io_VwirePorts_1_0_13_in( ArrayRowModule_1_io_V_wire_out_13 ),
       .io_VwirePorts_1_0_13_en( T381 ),
       .io_VwirePorts_1_0_13_out( VwireModule_io_VwirePorts_1_0_13_out ),
       .io_VwirePorts_1_0_12_in( ArrayRowModule_1_io_V_wire_out_12 ),
       .io_VwirePorts_1_0_12_en( T380 ),
       .io_VwirePorts_1_0_12_out( VwireModule_io_VwirePorts_1_0_12_out ),
       .io_VwirePorts_1_0_11_in( ArrayRowModule_1_io_V_wire_out_11 ),
       .io_VwirePorts_1_0_11_en( T379 ),
       .io_VwirePorts_1_0_11_out( VwireModule_io_VwirePorts_1_0_11_out ),
       .io_VwirePorts_1_0_10_in( ArrayRowModule_1_io_V_wire_out_10 ),
       .io_VwirePorts_1_0_10_en( T378 ),
       .io_VwirePorts_1_0_10_out( VwireModule_io_VwirePorts_1_0_10_out ),
       .io_VwirePorts_1_0_9_in( ArrayRowModule_1_io_V_wire_out_9 ),
       .io_VwirePorts_1_0_9_en( T377 ),
       .io_VwirePorts_1_0_9_out( VwireModule_io_VwirePorts_1_0_9_out ),
       .io_VwirePorts_1_0_8_in( ArrayRowModule_1_io_V_wire_out_8 ),
       .io_VwirePorts_1_0_8_en( T376 ),
       .io_VwirePorts_1_0_8_out( VwireModule_io_VwirePorts_1_0_8_out ),
       .io_VwirePorts_1_0_7_in( ArrayRowModule_1_io_V_wire_out_7 ),
       .io_VwirePorts_1_0_7_en( T375 ),
       .io_VwirePorts_1_0_7_out( VwireModule_io_VwirePorts_1_0_7_out ),
       .io_VwirePorts_1_0_6_in( ArrayRowModule_1_io_V_wire_out_6 ),
       .io_VwirePorts_1_0_6_en( T374 ),
       .io_VwirePorts_1_0_6_out( VwireModule_io_VwirePorts_1_0_6_out ),
       .io_VwirePorts_1_0_5_in( ArrayRowModule_1_io_V_wire_out_5 ),
       .io_VwirePorts_1_0_5_en( T373 ),
       .io_VwirePorts_1_0_5_out( VwireModule_io_VwirePorts_1_0_5_out ),
       .io_VwirePorts_1_0_4_in( ArrayRowModule_1_io_V_wire_out_4 ),
       .io_VwirePorts_1_0_4_en( T372 ),
       .io_VwirePorts_1_0_4_out( VwireModule_io_VwirePorts_1_0_4_out ),
       .io_VwirePorts_1_0_3_in( ArrayRowModule_1_io_V_wire_out_3 ),
       .io_VwirePorts_1_0_3_en( T371 ),
       .io_VwirePorts_1_0_3_out( VwireModule_io_VwirePorts_1_0_3_out ),
       .io_VwirePorts_1_0_2_in( ArrayRowModule_1_io_V_wire_out_2 ),
       .io_VwirePorts_1_0_2_en( T370 ),
       .io_VwirePorts_1_0_2_out( VwireModule_io_VwirePorts_1_0_2_out ),
       .io_VwirePorts_1_0_1_in( ArrayRowModule_1_io_V_wire_out_1 ),
       .io_VwirePorts_1_0_1_en( T369 ),
       .io_VwirePorts_1_0_1_out( VwireModule_io_VwirePorts_1_0_1_out ),
       .io_VwirePorts_1_0_0_in( ArrayRowModule_1_io_V_wire_out_0 ),
       .io_VwirePorts_1_0_0_en( T368 ),
       .io_VwirePorts_1_0_0_out( VwireModule_io_VwirePorts_1_0_0_out ),
       .io_VwirePorts_0_22_15_in( ArrayRowModule_io_V_wire_out_367 ),
       .io_VwirePorts_0_22_15_en( T367 ),
       .io_VwirePorts_0_22_15_out( VwireModule_io_VwirePorts_0_22_15_out ),
       .io_VwirePorts_0_22_14_in( ArrayRowModule_io_V_wire_out_366 ),
       .io_VwirePorts_0_22_14_en( T366 ),
       .io_VwirePorts_0_22_14_out( VwireModule_io_VwirePorts_0_22_14_out ),
       .io_VwirePorts_0_22_13_in( ArrayRowModule_io_V_wire_out_365 ),
       .io_VwirePorts_0_22_13_en( T365 ),
       .io_VwirePorts_0_22_13_out( VwireModule_io_VwirePorts_0_22_13_out ),
       .io_VwirePorts_0_22_12_in( ArrayRowModule_io_V_wire_out_364 ),
       .io_VwirePorts_0_22_12_en( T364 ),
       .io_VwirePorts_0_22_12_out( VwireModule_io_VwirePorts_0_22_12_out ),
       .io_VwirePorts_0_22_11_in( ArrayRowModule_io_V_wire_out_363 ),
       .io_VwirePorts_0_22_11_en( T363 ),
       .io_VwirePorts_0_22_11_out( VwireModule_io_VwirePorts_0_22_11_out ),
       .io_VwirePorts_0_22_10_in( ArrayRowModule_io_V_wire_out_362 ),
       .io_VwirePorts_0_22_10_en( T362 ),
       .io_VwirePorts_0_22_10_out( VwireModule_io_VwirePorts_0_22_10_out ),
       .io_VwirePorts_0_22_9_in( ArrayRowModule_io_V_wire_out_361 ),
       .io_VwirePorts_0_22_9_en( T361 ),
       .io_VwirePorts_0_22_9_out( VwireModule_io_VwirePorts_0_22_9_out ),
       .io_VwirePorts_0_22_8_in( ArrayRowModule_io_V_wire_out_360 ),
       .io_VwirePorts_0_22_8_en( T360 ),
       .io_VwirePorts_0_22_8_out( VwireModule_io_VwirePorts_0_22_8_out ),
       .io_VwirePorts_0_22_7_in( ArrayRowModule_io_V_wire_out_359 ),
       .io_VwirePorts_0_22_7_en( T359 ),
       .io_VwirePorts_0_22_7_out( VwireModule_io_VwirePorts_0_22_7_out ),
       .io_VwirePorts_0_22_6_in( ArrayRowModule_io_V_wire_out_358 ),
       .io_VwirePorts_0_22_6_en( T358 ),
       .io_VwirePorts_0_22_6_out( VwireModule_io_VwirePorts_0_22_6_out ),
       .io_VwirePorts_0_22_5_in( ArrayRowModule_io_V_wire_out_357 ),
       .io_VwirePorts_0_22_5_en( T357 ),
       .io_VwirePorts_0_22_5_out( VwireModule_io_VwirePorts_0_22_5_out ),
       .io_VwirePorts_0_22_4_in( ArrayRowModule_io_V_wire_out_356 ),
       .io_VwirePorts_0_22_4_en( T356 ),
       .io_VwirePorts_0_22_4_out( VwireModule_io_VwirePorts_0_22_4_out ),
       .io_VwirePorts_0_22_3_in( ArrayRowModule_io_V_wire_out_355 ),
       .io_VwirePorts_0_22_3_en( T355 ),
       .io_VwirePorts_0_22_3_out( VwireModule_io_VwirePorts_0_22_3_out ),
       .io_VwirePorts_0_22_2_in( ArrayRowModule_io_V_wire_out_354 ),
       .io_VwirePorts_0_22_2_en( T354 ),
       .io_VwirePorts_0_22_2_out( VwireModule_io_VwirePorts_0_22_2_out ),
       .io_VwirePorts_0_22_1_in( ArrayRowModule_io_V_wire_out_353 ),
       .io_VwirePorts_0_22_1_en( T353 ),
       .io_VwirePorts_0_22_1_out( VwireModule_io_VwirePorts_0_22_1_out ),
       .io_VwirePorts_0_22_0_in( ArrayRowModule_io_V_wire_out_352 ),
       .io_VwirePorts_0_22_0_en( T352 ),
       .io_VwirePorts_0_22_0_out( VwireModule_io_VwirePorts_0_22_0_out ),
       .io_VwirePorts_0_21_15_in( ArrayRowModule_io_V_wire_out_351 ),
       .io_VwirePorts_0_21_15_en( T351 ),
       .io_VwirePorts_0_21_15_out( VwireModule_io_VwirePorts_0_21_15_out ),
       .io_VwirePorts_0_21_14_in( ArrayRowModule_io_V_wire_out_350 ),
       .io_VwirePorts_0_21_14_en( T350 ),
       .io_VwirePorts_0_21_14_out( VwireModule_io_VwirePorts_0_21_14_out ),
       .io_VwirePorts_0_21_13_in( ArrayRowModule_io_V_wire_out_349 ),
       .io_VwirePorts_0_21_13_en( T349 ),
       .io_VwirePorts_0_21_13_out( VwireModule_io_VwirePorts_0_21_13_out ),
       .io_VwirePorts_0_21_12_in( ArrayRowModule_io_V_wire_out_348 ),
       .io_VwirePorts_0_21_12_en( T348 ),
       .io_VwirePorts_0_21_12_out( VwireModule_io_VwirePorts_0_21_12_out ),
       .io_VwirePorts_0_21_11_in( ArrayRowModule_io_V_wire_out_347 ),
       .io_VwirePorts_0_21_11_en( T347 ),
       .io_VwirePorts_0_21_11_out( VwireModule_io_VwirePorts_0_21_11_out ),
       .io_VwirePorts_0_21_10_in( ArrayRowModule_io_V_wire_out_346 ),
       .io_VwirePorts_0_21_10_en( T346 ),
       .io_VwirePorts_0_21_10_out( VwireModule_io_VwirePorts_0_21_10_out ),
       .io_VwirePorts_0_21_9_in( ArrayRowModule_io_V_wire_out_345 ),
       .io_VwirePorts_0_21_9_en( T345 ),
       .io_VwirePorts_0_21_9_out( VwireModule_io_VwirePorts_0_21_9_out ),
       .io_VwirePorts_0_21_8_in( ArrayRowModule_io_V_wire_out_344 ),
       .io_VwirePorts_0_21_8_en( T344 ),
       .io_VwirePorts_0_21_8_out( VwireModule_io_VwirePorts_0_21_8_out ),
       .io_VwirePorts_0_21_7_in( ArrayRowModule_io_V_wire_out_343 ),
       .io_VwirePorts_0_21_7_en( T343 ),
       .io_VwirePorts_0_21_7_out( VwireModule_io_VwirePorts_0_21_7_out ),
       .io_VwirePorts_0_21_6_in( ArrayRowModule_io_V_wire_out_342 ),
       .io_VwirePorts_0_21_6_en( T342 ),
       .io_VwirePorts_0_21_6_out( VwireModule_io_VwirePorts_0_21_6_out ),
       .io_VwirePorts_0_21_5_in( ArrayRowModule_io_V_wire_out_341 ),
       .io_VwirePorts_0_21_5_en( T341 ),
       .io_VwirePorts_0_21_5_out( VwireModule_io_VwirePorts_0_21_5_out ),
       .io_VwirePorts_0_21_4_in( ArrayRowModule_io_V_wire_out_340 ),
       .io_VwirePorts_0_21_4_en( T340 ),
       .io_VwirePorts_0_21_4_out( VwireModule_io_VwirePorts_0_21_4_out ),
       .io_VwirePorts_0_21_3_in( ArrayRowModule_io_V_wire_out_339 ),
       .io_VwirePorts_0_21_3_en( T339 ),
       .io_VwirePorts_0_21_3_out( VwireModule_io_VwirePorts_0_21_3_out ),
       .io_VwirePorts_0_21_2_in( ArrayRowModule_io_V_wire_out_338 ),
       .io_VwirePorts_0_21_2_en( T338 ),
       .io_VwirePorts_0_21_2_out( VwireModule_io_VwirePorts_0_21_2_out ),
       .io_VwirePorts_0_21_1_in( ArrayRowModule_io_V_wire_out_337 ),
       .io_VwirePorts_0_21_1_en( T337 ),
       .io_VwirePorts_0_21_1_out( VwireModule_io_VwirePorts_0_21_1_out ),
       .io_VwirePorts_0_21_0_in( ArrayRowModule_io_V_wire_out_336 ),
       .io_VwirePorts_0_21_0_en( T336 ),
       .io_VwirePorts_0_21_0_out( VwireModule_io_VwirePorts_0_21_0_out ),
       .io_VwirePorts_0_20_15_in( ArrayRowModule_io_V_wire_out_335 ),
       .io_VwirePorts_0_20_15_en( T335 ),
       .io_VwirePorts_0_20_15_out( VwireModule_io_VwirePorts_0_20_15_out ),
       .io_VwirePorts_0_20_14_in( ArrayRowModule_io_V_wire_out_334 ),
       .io_VwirePorts_0_20_14_en( T334 ),
       .io_VwirePorts_0_20_14_out( VwireModule_io_VwirePorts_0_20_14_out ),
       .io_VwirePorts_0_20_13_in( ArrayRowModule_io_V_wire_out_333 ),
       .io_VwirePorts_0_20_13_en( T333 ),
       .io_VwirePorts_0_20_13_out( VwireModule_io_VwirePorts_0_20_13_out ),
       .io_VwirePorts_0_20_12_in( ArrayRowModule_io_V_wire_out_332 ),
       .io_VwirePorts_0_20_12_en( T332 ),
       .io_VwirePorts_0_20_12_out( VwireModule_io_VwirePorts_0_20_12_out ),
       .io_VwirePorts_0_20_11_in( ArrayRowModule_io_V_wire_out_331 ),
       .io_VwirePorts_0_20_11_en( T331 ),
       .io_VwirePorts_0_20_11_out( VwireModule_io_VwirePorts_0_20_11_out ),
       .io_VwirePorts_0_20_10_in( ArrayRowModule_io_V_wire_out_330 ),
       .io_VwirePorts_0_20_10_en( T330 ),
       .io_VwirePorts_0_20_10_out( VwireModule_io_VwirePorts_0_20_10_out ),
       .io_VwirePorts_0_20_9_in( ArrayRowModule_io_V_wire_out_329 ),
       .io_VwirePorts_0_20_9_en( T329 ),
       .io_VwirePorts_0_20_9_out( VwireModule_io_VwirePorts_0_20_9_out ),
       .io_VwirePorts_0_20_8_in( ArrayRowModule_io_V_wire_out_328 ),
       .io_VwirePorts_0_20_8_en( T328 ),
       .io_VwirePorts_0_20_8_out( VwireModule_io_VwirePorts_0_20_8_out ),
       .io_VwirePorts_0_20_7_in( ArrayRowModule_io_V_wire_out_327 ),
       .io_VwirePorts_0_20_7_en( T327 ),
       .io_VwirePorts_0_20_7_out( VwireModule_io_VwirePorts_0_20_7_out ),
       .io_VwirePorts_0_20_6_in( ArrayRowModule_io_V_wire_out_326 ),
       .io_VwirePorts_0_20_6_en( T326 ),
       .io_VwirePorts_0_20_6_out( VwireModule_io_VwirePorts_0_20_6_out ),
       .io_VwirePorts_0_20_5_in( ArrayRowModule_io_V_wire_out_325 ),
       .io_VwirePorts_0_20_5_en( T325 ),
       .io_VwirePorts_0_20_5_out( VwireModule_io_VwirePorts_0_20_5_out ),
       .io_VwirePorts_0_20_4_in( ArrayRowModule_io_V_wire_out_324 ),
       .io_VwirePorts_0_20_4_en( T324 ),
       .io_VwirePorts_0_20_4_out( VwireModule_io_VwirePorts_0_20_4_out ),
       .io_VwirePorts_0_20_3_in( ArrayRowModule_io_V_wire_out_323 ),
       .io_VwirePorts_0_20_3_en( T323 ),
       .io_VwirePorts_0_20_3_out( VwireModule_io_VwirePorts_0_20_3_out ),
       .io_VwirePorts_0_20_2_in( ArrayRowModule_io_V_wire_out_322 ),
       .io_VwirePorts_0_20_2_en( T322 ),
       .io_VwirePorts_0_20_2_out( VwireModule_io_VwirePorts_0_20_2_out ),
       .io_VwirePorts_0_20_1_in( ArrayRowModule_io_V_wire_out_321 ),
       .io_VwirePorts_0_20_1_en( T321 ),
       .io_VwirePorts_0_20_1_out( VwireModule_io_VwirePorts_0_20_1_out ),
       .io_VwirePorts_0_20_0_in( ArrayRowModule_io_V_wire_out_320 ),
       .io_VwirePorts_0_20_0_en( T320 ),
       .io_VwirePorts_0_20_0_out( VwireModule_io_VwirePorts_0_20_0_out ),
       .io_VwirePorts_0_19_15_in( ArrayRowModule_io_V_wire_out_319 ),
       .io_VwirePorts_0_19_15_en( T319 ),
       .io_VwirePorts_0_19_15_out( VwireModule_io_VwirePorts_0_19_15_out ),
       .io_VwirePorts_0_19_14_in( ArrayRowModule_io_V_wire_out_318 ),
       .io_VwirePorts_0_19_14_en( T318 ),
       .io_VwirePorts_0_19_14_out( VwireModule_io_VwirePorts_0_19_14_out ),
       .io_VwirePorts_0_19_13_in( ArrayRowModule_io_V_wire_out_317 ),
       .io_VwirePorts_0_19_13_en( T317 ),
       .io_VwirePorts_0_19_13_out( VwireModule_io_VwirePorts_0_19_13_out ),
       .io_VwirePorts_0_19_12_in( ArrayRowModule_io_V_wire_out_316 ),
       .io_VwirePorts_0_19_12_en( T316 ),
       .io_VwirePorts_0_19_12_out( VwireModule_io_VwirePorts_0_19_12_out ),
       .io_VwirePorts_0_19_11_in( ArrayRowModule_io_V_wire_out_315 ),
       .io_VwirePorts_0_19_11_en( T315 ),
       .io_VwirePorts_0_19_11_out( VwireModule_io_VwirePorts_0_19_11_out ),
       .io_VwirePorts_0_19_10_in( ArrayRowModule_io_V_wire_out_314 ),
       .io_VwirePorts_0_19_10_en( T314 ),
       .io_VwirePorts_0_19_10_out( VwireModule_io_VwirePorts_0_19_10_out ),
       .io_VwirePorts_0_19_9_in( ArrayRowModule_io_V_wire_out_313 ),
       .io_VwirePorts_0_19_9_en( T313 ),
       .io_VwirePorts_0_19_9_out( VwireModule_io_VwirePorts_0_19_9_out ),
       .io_VwirePorts_0_19_8_in( ArrayRowModule_io_V_wire_out_312 ),
       .io_VwirePorts_0_19_8_en( T312 ),
       .io_VwirePorts_0_19_8_out( VwireModule_io_VwirePorts_0_19_8_out ),
       .io_VwirePorts_0_19_7_in( ArrayRowModule_io_V_wire_out_311 ),
       .io_VwirePorts_0_19_7_en( T311 ),
       .io_VwirePorts_0_19_7_out( VwireModule_io_VwirePorts_0_19_7_out ),
       .io_VwirePorts_0_19_6_in( ArrayRowModule_io_V_wire_out_310 ),
       .io_VwirePorts_0_19_6_en( T310 ),
       .io_VwirePorts_0_19_6_out( VwireModule_io_VwirePorts_0_19_6_out ),
       .io_VwirePorts_0_19_5_in( ArrayRowModule_io_V_wire_out_309 ),
       .io_VwirePorts_0_19_5_en( T309 ),
       .io_VwirePorts_0_19_5_out( VwireModule_io_VwirePorts_0_19_5_out ),
       .io_VwirePorts_0_19_4_in( ArrayRowModule_io_V_wire_out_308 ),
       .io_VwirePorts_0_19_4_en( T308 ),
       .io_VwirePorts_0_19_4_out( VwireModule_io_VwirePorts_0_19_4_out ),
       .io_VwirePorts_0_19_3_in( ArrayRowModule_io_V_wire_out_307 ),
       .io_VwirePorts_0_19_3_en( T307 ),
       .io_VwirePorts_0_19_3_out( VwireModule_io_VwirePorts_0_19_3_out ),
       .io_VwirePorts_0_19_2_in( ArrayRowModule_io_V_wire_out_306 ),
       .io_VwirePorts_0_19_2_en( T306 ),
       .io_VwirePorts_0_19_2_out( VwireModule_io_VwirePorts_0_19_2_out ),
       .io_VwirePorts_0_19_1_in( ArrayRowModule_io_V_wire_out_305 ),
       .io_VwirePorts_0_19_1_en( T305 ),
       .io_VwirePorts_0_19_1_out( VwireModule_io_VwirePorts_0_19_1_out ),
       .io_VwirePorts_0_19_0_in( ArrayRowModule_io_V_wire_out_304 ),
       .io_VwirePorts_0_19_0_en( T304 ),
       .io_VwirePorts_0_19_0_out( VwireModule_io_VwirePorts_0_19_0_out ),
       .io_VwirePorts_0_18_15_in( ArrayRowModule_io_V_wire_out_303 ),
       .io_VwirePorts_0_18_15_en( T303 ),
       .io_VwirePorts_0_18_15_out( VwireModule_io_VwirePorts_0_18_15_out ),
       .io_VwirePorts_0_18_14_in( ArrayRowModule_io_V_wire_out_302 ),
       .io_VwirePorts_0_18_14_en( T302 ),
       .io_VwirePorts_0_18_14_out( VwireModule_io_VwirePorts_0_18_14_out ),
       .io_VwirePorts_0_18_13_in( ArrayRowModule_io_V_wire_out_301 ),
       .io_VwirePorts_0_18_13_en( T301 ),
       .io_VwirePorts_0_18_13_out( VwireModule_io_VwirePorts_0_18_13_out ),
       .io_VwirePorts_0_18_12_in( ArrayRowModule_io_V_wire_out_300 ),
       .io_VwirePorts_0_18_12_en( T300 ),
       .io_VwirePorts_0_18_12_out( VwireModule_io_VwirePorts_0_18_12_out ),
       .io_VwirePorts_0_18_11_in( ArrayRowModule_io_V_wire_out_299 ),
       .io_VwirePorts_0_18_11_en( T299 ),
       .io_VwirePorts_0_18_11_out( VwireModule_io_VwirePorts_0_18_11_out ),
       .io_VwirePorts_0_18_10_in( ArrayRowModule_io_V_wire_out_298 ),
       .io_VwirePorts_0_18_10_en( T298 ),
       .io_VwirePorts_0_18_10_out( VwireModule_io_VwirePorts_0_18_10_out ),
       .io_VwirePorts_0_18_9_in( ArrayRowModule_io_V_wire_out_297 ),
       .io_VwirePorts_0_18_9_en( T297 ),
       .io_VwirePorts_0_18_9_out( VwireModule_io_VwirePorts_0_18_9_out ),
       .io_VwirePorts_0_18_8_in( ArrayRowModule_io_V_wire_out_296 ),
       .io_VwirePorts_0_18_8_en( T296 ),
       .io_VwirePorts_0_18_8_out( VwireModule_io_VwirePorts_0_18_8_out ),
       .io_VwirePorts_0_18_7_in( ArrayRowModule_io_V_wire_out_295 ),
       .io_VwirePorts_0_18_7_en( T295 ),
       .io_VwirePorts_0_18_7_out( VwireModule_io_VwirePorts_0_18_7_out ),
       .io_VwirePorts_0_18_6_in( ArrayRowModule_io_V_wire_out_294 ),
       .io_VwirePorts_0_18_6_en( T294 ),
       .io_VwirePorts_0_18_6_out( VwireModule_io_VwirePorts_0_18_6_out ),
       .io_VwirePorts_0_18_5_in( ArrayRowModule_io_V_wire_out_293 ),
       .io_VwirePorts_0_18_5_en( T293 ),
       .io_VwirePorts_0_18_5_out( VwireModule_io_VwirePorts_0_18_5_out ),
       .io_VwirePorts_0_18_4_in( ArrayRowModule_io_V_wire_out_292 ),
       .io_VwirePorts_0_18_4_en( T292 ),
       .io_VwirePorts_0_18_4_out( VwireModule_io_VwirePorts_0_18_4_out ),
       .io_VwirePorts_0_18_3_in( ArrayRowModule_io_V_wire_out_291 ),
       .io_VwirePorts_0_18_3_en( T291 ),
       .io_VwirePorts_0_18_3_out( VwireModule_io_VwirePorts_0_18_3_out ),
       .io_VwirePorts_0_18_2_in( ArrayRowModule_io_V_wire_out_290 ),
       .io_VwirePorts_0_18_2_en( T290 ),
       .io_VwirePorts_0_18_2_out( VwireModule_io_VwirePorts_0_18_2_out ),
       .io_VwirePorts_0_18_1_in( ArrayRowModule_io_V_wire_out_289 ),
       .io_VwirePorts_0_18_1_en( T289 ),
       .io_VwirePorts_0_18_1_out( VwireModule_io_VwirePorts_0_18_1_out ),
       .io_VwirePorts_0_18_0_in( ArrayRowModule_io_V_wire_out_288 ),
       .io_VwirePorts_0_18_0_en( T288 ),
       .io_VwirePorts_0_18_0_out( VwireModule_io_VwirePorts_0_18_0_out ),
       .io_VwirePorts_0_17_15_in( ArrayRowModule_io_V_wire_out_287 ),
       .io_VwirePorts_0_17_15_en( T287 ),
       .io_VwirePorts_0_17_15_out( VwireModule_io_VwirePorts_0_17_15_out ),
       .io_VwirePorts_0_17_14_in( ArrayRowModule_io_V_wire_out_286 ),
       .io_VwirePorts_0_17_14_en( T286 ),
       .io_VwirePorts_0_17_14_out( VwireModule_io_VwirePorts_0_17_14_out ),
       .io_VwirePorts_0_17_13_in( ArrayRowModule_io_V_wire_out_285 ),
       .io_VwirePorts_0_17_13_en( T285 ),
       .io_VwirePorts_0_17_13_out( VwireModule_io_VwirePorts_0_17_13_out ),
       .io_VwirePorts_0_17_12_in( ArrayRowModule_io_V_wire_out_284 ),
       .io_VwirePorts_0_17_12_en( T284 ),
       .io_VwirePorts_0_17_12_out( VwireModule_io_VwirePorts_0_17_12_out ),
       .io_VwirePorts_0_17_11_in( ArrayRowModule_io_V_wire_out_283 ),
       .io_VwirePorts_0_17_11_en( T283 ),
       .io_VwirePorts_0_17_11_out( VwireModule_io_VwirePorts_0_17_11_out ),
       .io_VwirePorts_0_17_10_in( ArrayRowModule_io_V_wire_out_282 ),
       .io_VwirePorts_0_17_10_en( T282 ),
       .io_VwirePorts_0_17_10_out( VwireModule_io_VwirePorts_0_17_10_out ),
       .io_VwirePorts_0_17_9_in( ArrayRowModule_io_V_wire_out_281 ),
       .io_VwirePorts_0_17_9_en( T281 ),
       .io_VwirePorts_0_17_9_out( VwireModule_io_VwirePorts_0_17_9_out ),
       .io_VwirePorts_0_17_8_in( ArrayRowModule_io_V_wire_out_280 ),
       .io_VwirePorts_0_17_8_en( T280 ),
       .io_VwirePorts_0_17_8_out( VwireModule_io_VwirePorts_0_17_8_out ),
       .io_VwirePorts_0_17_7_in( ArrayRowModule_io_V_wire_out_279 ),
       .io_VwirePorts_0_17_7_en( T279 ),
       .io_VwirePorts_0_17_7_out( VwireModule_io_VwirePorts_0_17_7_out ),
       .io_VwirePorts_0_17_6_in( ArrayRowModule_io_V_wire_out_278 ),
       .io_VwirePorts_0_17_6_en( T278 ),
       .io_VwirePorts_0_17_6_out( VwireModule_io_VwirePorts_0_17_6_out ),
       .io_VwirePorts_0_17_5_in( ArrayRowModule_io_V_wire_out_277 ),
       .io_VwirePorts_0_17_5_en( T277 ),
       .io_VwirePorts_0_17_5_out( VwireModule_io_VwirePorts_0_17_5_out ),
       .io_VwirePorts_0_17_4_in( ArrayRowModule_io_V_wire_out_276 ),
       .io_VwirePorts_0_17_4_en( T276 ),
       .io_VwirePorts_0_17_4_out( VwireModule_io_VwirePorts_0_17_4_out ),
       .io_VwirePorts_0_17_3_in( ArrayRowModule_io_V_wire_out_275 ),
       .io_VwirePorts_0_17_3_en( T275 ),
       .io_VwirePorts_0_17_3_out( VwireModule_io_VwirePorts_0_17_3_out ),
       .io_VwirePorts_0_17_2_in( ArrayRowModule_io_V_wire_out_274 ),
       .io_VwirePorts_0_17_2_en( T274 ),
       .io_VwirePorts_0_17_2_out( VwireModule_io_VwirePorts_0_17_2_out ),
       .io_VwirePorts_0_17_1_in( ArrayRowModule_io_V_wire_out_273 ),
       .io_VwirePorts_0_17_1_en( T273 ),
       .io_VwirePorts_0_17_1_out( VwireModule_io_VwirePorts_0_17_1_out ),
       .io_VwirePorts_0_17_0_in( ArrayRowModule_io_V_wire_out_272 ),
       .io_VwirePorts_0_17_0_en( T272 ),
       .io_VwirePorts_0_17_0_out( VwireModule_io_VwirePorts_0_17_0_out ),
       .io_VwirePorts_0_16_15_in( ArrayRowModule_io_V_wire_out_271 ),
       .io_VwirePorts_0_16_15_en( T271 ),
       .io_VwirePorts_0_16_15_out( VwireModule_io_VwirePorts_0_16_15_out ),
       .io_VwirePorts_0_16_14_in( ArrayRowModule_io_V_wire_out_270 ),
       .io_VwirePorts_0_16_14_en( T270 ),
       .io_VwirePorts_0_16_14_out( VwireModule_io_VwirePorts_0_16_14_out ),
       .io_VwirePorts_0_16_13_in( ArrayRowModule_io_V_wire_out_269 ),
       .io_VwirePorts_0_16_13_en( T269 ),
       .io_VwirePorts_0_16_13_out( VwireModule_io_VwirePorts_0_16_13_out ),
       .io_VwirePorts_0_16_12_in( ArrayRowModule_io_V_wire_out_268 ),
       .io_VwirePorts_0_16_12_en( T268 ),
       .io_VwirePorts_0_16_12_out( VwireModule_io_VwirePorts_0_16_12_out ),
       .io_VwirePorts_0_16_11_in( ArrayRowModule_io_V_wire_out_267 ),
       .io_VwirePorts_0_16_11_en( T267 ),
       .io_VwirePorts_0_16_11_out( VwireModule_io_VwirePorts_0_16_11_out ),
       .io_VwirePorts_0_16_10_in( ArrayRowModule_io_V_wire_out_266 ),
       .io_VwirePorts_0_16_10_en( T266 ),
       .io_VwirePorts_0_16_10_out( VwireModule_io_VwirePorts_0_16_10_out ),
       .io_VwirePorts_0_16_9_in( ArrayRowModule_io_V_wire_out_265 ),
       .io_VwirePorts_0_16_9_en( T265 ),
       .io_VwirePorts_0_16_9_out( VwireModule_io_VwirePorts_0_16_9_out ),
       .io_VwirePorts_0_16_8_in( ArrayRowModule_io_V_wire_out_264 ),
       .io_VwirePorts_0_16_8_en( T264 ),
       .io_VwirePorts_0_16_8_out( VwireModule_io_VwirePorts_0_16_8_out ),
       .io_VwirePorts_0_16_7_in( ArrayRowModule_io_V_wire_out_263 ),
       .io_VwirePorts_0_16_7_en( T263 ),
       .io_VwirePorts_0_16_7_out( VwireModule_io_VwirePorts_0_16_7_out ),
       .io_VwirePorts_0_16_6_in( ArrayRowModule_io_V_wire_out_262 ),
       .io_VwirePorts_0_16_6_en( T262 ),
       .io_VwirePorts_0_16_6_out( VwireModule_io_VwirePorts_0_16_6_out ),
       .io_VwirePorts_0_16_5_in( ArrayRowModule_io_V_wire_out_261 ),
       .io_VwirePorts_0_16_5_en( T261 ),
       .io_VwirePorts_0_16_5_out( VwireModule_io_VwirePorts_0_16_5_out ),
       .io_VwirePorts_0_16_4_in( ArrayRowModule_io_V_wire_out_260 ),
       .io_VwirePorts_0_16_4_en( T260 ),
       .io_VwirePorts_0_16_4_out( VwireModule_io_VwirePorts_0_16_4_out ),
       .io_VwirePorts_0_16_3_in( ArrayRowModule_io_V_wire_out_259 ),
       .io_VwirePorts_0_16_3_en( T259 ),
       .io_VwirePorts_0_16_3_out( VwireModule_io_VwirePorts_0_16_3_out ),
       .io_VwirePorts_0_16_2_in( ArrayRowModule_io_V_wire_out_258 ),
       .io_VwirePorts_0_16_2_en( T258 ),
       .io_VwirePorts_0_16_2_out( VwireModule_io_VwirePorts_0_16_2_out ),
       .io_VwirePorts_0_16_1_in( ArrayRowModule_io_V_wire_out_257 ),
       .io_VwirePorts_0_16_1_en( T257 ),
       .io_VwirePorts_0_16_1_out( VwireModule_io_VwirePorts_0_16_1_out ),
       .io_VwirePorts_0_16_0_in( ArrayRowModule_io_V_wire_out_256 ),
       .io_VwirePorts_0_16_0_en( T256 ),
       .io_VwirePorts_0_16_0_out( VwireModule_io_VwirePorts_0_16_0_out ),
       .io_VwirePorts_0_15_15_in( ArrayRowModule_io_V_wire_out_255 ),
       .io_VwirePorts_0_15_15_en( T255 ),
       .io_VwirePorts_0_15_15_out( VwireModule_io_VwirePorts_0_15_15_out ),
       .io_VwirePorts_0_15_14_in( ArrayRowModule_io_V_wire_out_254 ),
       .io_VwirePorts_0_15_14_en( T254 ),
       .io_VwirePorts_0_15_14_out( VwireModule_io_VwirePorts_0_15_14_out ),
       .io_VwirePorts_0_15_13_in( ArrayRowModule_io_V_wire_out_253 ),
       .io_VwirePorts_0_15_13_en( T253 ),
       .io_VwirePorts_0_15_13_out( VwireModule_io_VwirePorts_0_15_13_out ),
       .io_VwirePorts_0_15_12_in( ArrayRowModule_io_V_wire_out_252 ),
       .io_VwirePorts_0_15_12_en( T252 ),
       .io_VwirePorts_0_15_12_out( VwireModule_io_VwirePorts_0_15_12_out ),
       .io_VwirePorts_0_15_11_in( ArrayRowModule_io_V_wire_out_251 ),
       .io_VwirePorts_0_15_11_en( T251 ),
       .io_VwirePorts_0_15_11_out( VwireModule_io_VwirePorts_0_15_11_out ),
       .io_VwirePorts_0_15_10_in( ArrayRowModule_io_V_wire_out_250 ),
       .io_VwirePorts_0_15_10_en( T250 ),
       .io_VwirePorts_0_15_10_out( VwireModule_io_VwirePorts_0_15_10_out ),
       .io_VwirePorts_0_15_9_in( ArrayRowModule_io_V_wire_out_249 ),
       .io_VwirePorts_0_15_9_en( T249 ),
       .io_VwirePorts_0_15_9_out( VwireModule_io_VwirePorts_0_15_9_out ),
       .io_VwirePorts_0_15_8_in( ArrayRowModule_io_V_wire_out_248 ),
       .io_VwirePorts_0_15_8_en( T248 ),
       .io_VwirePorts_0_15_8_out( VwireModule_io_VwirePorts_0_15_8_out ),
       .io_VwirePorts_0_15_7_in( ArrayRowModule_io_V_wire_out_247 ),
       .io_VwirePorts_0_15_7_en( T247 ),
       .io_VwirePorts_0_15_7_out( VwireModule_io_VwirePorts_0_15_7_out ),
       .io_VwirePorts_0_15_6_in( ArrayRowModule_io_V_wire_out_246 ),
       .io_VwirePorts_0_15_6_en( T246 ),
       .io_VwirePorts_0_15_6_out( VwireModule_io_VwirePorts_0_15_6_out ),
       .io_VwirePorts_0_15_5_in( ArrayRowModule_io_V_wire_out_245 ),
       .io_VwirePorts_0_15_5_en( T245 ),
       .io_VwirePorts_0_15_5_out( VwireModule_io_VwirePorts_0_15_5_out ),
       .io_VwirePorts_0_15_4_in( ArrayRowModule_io_V_wire_out_244 ),
       .io_VwirePorts_0_15_4_en( T244 ),
       .io_VwirePorts_0_15_4_out( VwireModule_io_VwirePorts_0_15_4_out ),
       .io_VwirePorts_0_15_3_in( ArrayRowModule_io_V_wire_out_243 ),
       .io_VwirePorts_0_15_3_en( T243 ),
       .io_VwirePorts_0_15_3_out( VwireModule_io_VwirePorts_0_15_3_out ),
       .io_VwirePorts_0_15_2_in( ArrayRowModule_io_V_wire_out_242 ),
       .io_VwirePorts_0_15_2_en( T242 ),
       .io_VwirePorts_0_15_2_out( VwireModule_io_VwirePorts_0_15_2_out ),
       .io_VwirePorts_0_15_1_in( ArrayRowModule_io_V_wire_out_241 ),
       .io_VwirePorts_0_15_1_en( T241 ),
       .io_VwirePorts_0_15_1_out( VwireModule_io_VwirePorts_0_15_1_out ),
       .io_VwirePorts_0_15_0_in( ArrayRowModule_io_V_wire_out_240 ),
       .io_VwirePorts_0_15_0_en( T240 ),
       .io_VwirePorts_0_15_0_out( VwireModule_io_VwirePorts_0_15_0_out ),
       .io_VwirePorts_0_14_15_in( ArrayRowModule_io_V_wire_out_239 ),
       .io_VwirePorts_0_14_15_en( T239 ),
       .io_VwirePorts_0_14_15_out( VwireModule_io_VwirePorts_0_14_15_out ),
       .io_VwirePorts_0_14_14_in( ArrayRowModule_io_V_wire_out_238 ),
       .io_VwirePorts_0_14_14_en( T238 ),
       .io_VwirePorts_0_14_14_out( VwireModule_io_VwirePorts_0_14_14_out ),
       .io_VwirePorts_0_14_13_in( ArrayRowModule_io_V_wire_out_237 ),
       .io_VwirePorts_0_14_13_en( T237 ),
       .io_VwirePorts_0_14_13_out( VwireModule_io_VwirePorts_0_14_13_out ),
       .io_VwirePorts_0_14_12_in( ArrayRowModule_io_V_wire_out_236 ),
       .io_VwirePorts_0_14_12_en( T236 ),
       .io_VwirePorts_0_14_12_out( VwireModule_io_VwirePorts_0_14_12_out ),
       .io_VwirePorts_0_14_11_in( ArrayRowModule_io_V_wire_out_235 ),
       .io_VwirePorts_0_14_11_en( T235 ),
       .io_VwirePorts_0_14_11_out( VwireModule_io_VwirePorts_0_14_11_out ),
       .io_VwirePorts_0_14_10_in( ArrayRowModule_io_V_wire_out_234 ),
       .io_VwirePorts_0_14_10_en( T234 ),
       .io_VwirePorts_0_14_10_out( VwireModule_io_VwirePorts_0_14_10_out ),
       .io_VwirePorts_0_14_9_in( ArrayRowModule_io_V_wire_out_233 ),
       .io_VwirePorts_0_14_9_en( T233 ),
       .io_VwirePorts_0_14_9_out( VwireModule_io_VwirePorts_0_14_9_out ),
       .io_VwirePorts_0_14_8_in( ArrayRowModule_io_V_wire_out_232 ),
       .io_VwirePorts_0_14_8_en( T232 ),
       .io_VwirePorts_0_14_8_out( VwireModule_io_VwirePorts_0_14_8_out ),
       .io_VwirePorts_0_14_7_in( ArrayRowModule_io_V_wire_out_231 ),
       .io_VwirePorts_0_14_7_en( T231 ),
       .io_VwirePorts_0_14_7_out( VwireModule_io_VwirePorts_0_14_7_out ),
       .io_VwirePorts_0_14_6_in( ArrayRowModule_io_V_wire_out_230 ),
       .io_VwirePorts_0_14_6_en( T230 ),
       .io_VwirePorts_0_14_6_out( VwireModule_io_VwirePorts_0_14_6_out ),
       .io_VwirePorts_0_14_5_in( ArrayRowModule_io_V_wire_out_229 ),
       .io_VwirePorts_0_14_5_en( T229 ),
       .io_VwirePorts_0_14_5_out( VwireModule_io_VwirePorts_0_14_5_out ),
       .io_VwirePorts_0_14_4_in( ArrayRowModule_io_V_wire_out_228 ),
       .io_VwirePorts_0_14_4_en( T228 ),
       .io_VwirePorts_0_14_4_out( VwireModule_io_VwirePorts_0_14_4_out ),
       .io_VwirePorts_0_14_3_in( ArrayRowModule_io_V_wire_out_227 ),
       .io_VwirePorts_0_14_3_en( T227 ),
       .io_VwirePorts_0_14_3_out( VwireModule_io_VwirePorts_0_14_3_out ),
       .io_VwirePorts_0_14_2_in( ArrayRowModule_io_V_wire_out_226 ),
       .io_VwirePorts_0_14_2_en( T226 ),
       .io_VwirePorts_0_14_2_out( VwireModule_io_VwirePorts_0_14_2_out ),
       .io_VwirePorts_0_14_1_in( ArrayRowModule_io_V_wire_out_225 ),
       .io_VwirePorts_0_14_1_en( T225 ),
       .io_VwirePorts_0_14_1_out( VwireModule_io_VwirePorts_0_14_1_out ),
       .io_VwirePorts_0_14_0_in( ArrayRowModule_io_V_wire_out_224 ),
       .io_VwirePorts_0_14_0_en( T224 ),
       .io_VwirePorts_0_14_0_out( VwireModule_io_VwirePorts_0_14_0_out ),
       .io_VwirePorts_0_13_15_in( ArrayRowModule_io_V_wire_out_223 ),
       .io_VwirePorts_0_13_15_en( T223 ),
       .io_VwirePorts_0_13_15_out( VwireModule_io_VwirePorts_0_13_15_out ),
       .io_VwirePorts_0_13_14_in( ArrayRowModule_io_V_wire_out_222 ),
       .io_VwirePorts_0_13_14_en( T222 ),
       .io_VwirePorts_0_13_14_out( VwireModule_io_VwirePorts_0_13_14_out ),
       .io_VwirePorts_0_13_13_in( ArrayRowModule_io_V_wire_out_221 ),
       .io_VwirePorts_0_13_13_en( T221 ),
       .io_VwirePorts_0_13_13_out( VwireModule_io_VwirePorts_0_13_13_out ),
       .io_VwirePorts_0_13_12_in( ArrayRowModule_io_V_wire_out_220 ),
       .io_VwirePorts_0_13_12_en( T220 ),
       .io_VwirePorts_0_13_12_out( VwireModule_io_VwirePorts_0_13_12_out ),
       .io_VwirePorts_0_13_11_in( ArrayRowModule_io_V_wire_out_219 ),
       .io_VwirePorts_0_13_11_en( T219 ),
       .io_VwirePorts_0_13_11_out( VwireModule_io_VwirePorts_0_13_11_out ),
       .io_VwirePorts_0_13_10_in( ArrayRowModule_io_V_wire_out_218 ),
       .io_VwirePorts_0_13_10_en( T218 ),
       .io_VwirePorts_0_13_10_out( VwireModule_io_VwirePorts_0_13_10_out ),
       .io_VwirePorts_0_13_9_in( ArrayRowModule_io_V_wire_out_217 ),
       .io_VwirePorts_0_13_9_en( T217 ),
       .io_VwirePorts_0_13_9_out( VwireModule_io_VwirePorts_0_13_9_out ),
       .io_VwirePorts_0_13_8_in( ArrayRowModule_io_V_wire_out_216 ),
       .io_VwirePorts_0_13_8_en( T216 ),
       .io_VwirePorts_0_13_8_out( VwireModule_io_VwirePorts_0_13_8_out ),
       .io_VwirePorts_0_13_7_in( ArrayRowModule_io_V_wire_out_215 ),
       .io_VwirePorts_0_13_7_en( T215 ),
       .io_VwirePorts_0_13_7_out( VwireModule_io_VwirePorts_0_13_7_out ),
       .io_VwirePorts_0_13_6_in( ArrayRowModule_io_V_wire_out_214 ),
       .io_VwirePorts_0_13_6_en( T214 ),
       .io_VwirePorts_0_13_6_out( VwireModule_io_VwirePorts_0_13_6_out ),
       .io_VwirePorts_0_13_5_in( ArrayRowModule_io_V_wire_out_213 ),
       .io_VwirePorts_0_13_5_en( T213 ),
       .io_VwirePorts_0_13_5_out( VwireModule_io_VwirePorts_0_13_5_out ),
       .io_VwirePorts_0_13_4_in( ArrayRowModule_io_V_wire_out_212 ),
       .io_VwirePorts_0_13_4_en( T212 ),
       .io_VwirePorts_0_13_4_out( VwireModule_io_VwirePorts_0_13_4_out ),
       .io_VwirePorts_0_13_3_in( ArrayRowModule_io_V_wire_out_211 ),
       .io_VwirePorts_0_13_3_en( T211 ),
       .io_VwirePorts_0_13_3_out( VwireModule_io_VwirePorts_0_13_3_out ),
       .io_VwirePorts_0_13_2_in( ArrayRowModule_io_V_wire_out_210 ),
       .io_VwirePorts_0_13_2_en( T210 ),
       .io_VwirePorts_0_13_2_out( VwireModule_io_VwirePorts_0_13_2_out ),
       .io_VwirePorts_0_13_1_in( ArrayRowModule_io_V_wire_out_209 ),
       .io_VwirePorts_0_13_1_en( T209 ),
       .io_VwirePorts_0_13_1_out( VwireModule_io_VwirePorts_0_13_1_out ),
       .io_VwirePorts_0_13_0_in( ArrayRowModule_io_V_wire_out_208 ),
       .io_VwirePorts_0_13_0_en( T208 ),
       .io_VwirePorts_0_13_0_out( VwireModule_io_VwirePorts_0_13_0_out ),
       .io_VwirePorts_0_12_15_in( ArrayRowModule_io_V_wire_out_207 ),
       .io_VwirePorts_0_12_15_en( T207 ),
       .io_VwirePorts_0_12_15_out( VwireModule_io_VwirePorts_0_12_15_out ),
       .io_VwirePorts_0_12_14_in( ArrayRowModule_io_V_wire_out_206 ),
       .io_VwirePorts_0_12_14_en( T206 ),
       .io_VwirePorts_0_12_14_out( VwireModule_io_VwirePorts_0_12_14_out ),
       .io_VwirePorts_0_12_13_in( ArrayRowModule_io_V_wire_out_205 ),
       .io_VwirePorts_0_12_13_en( T205 ),
       .io_VwirePorts_0_12_13_out( VwireModule_io_VwirePorts_0_12_13_out ),
       .io_VwirePorts_0_12_12_in( ArrayRowModule_io_V_wire_out_204 ),
       .io_VwirePorts_0_12_12_en( T204 ),
       .io_VwirePorts_0_12_12_out( VwireModule_io_VwirePorts_0_12_12_out ),
       .io_VwirePorts_0_12_11_in( ArrayRowModule_io_V_wire_out_203 ),
       .io_VwirePorts_0_12_11_en( T203 ),
       .io_VwirePorts_0_12_11_out( VwireModule_io_VwirePorts_0_12_11_out ),
       .io_VwirePorts_0_12_10_in( ArrayRowModule_io_V_wire_out_202 ),
       .io_VwirePorts_0_12_10_en( T202 ),
       .io_VwirePorts_0_12_10_out( VwireModule_io_VwirePorts_0_12_10_out ),
       .io_VwirePorts_0_12_9_in( ArrayRowModule_io_V_wire_out_201 ),
       .io_VwirePorts_0_12_9_en( T201 ),
       .io_VwirePorts_0_12_9_out( VwireModule_io_VwirePorts_0_12_9_out ),
       .io_VwirePorts_0_12_8_in( ArrayRowModule_io_V_wire_out_200 ),
       .io_VwirePorts_0_12_8_en( T200 ),
       .io_VwirePorts_0_12_8_out( VwireModule_io_VwirePorts_0_12_8_out ),
       .io_VwirePorts_0_12_7_in( ArrayRowModule_io_V_wire_out_199 ),
       .io_VwirePorts_0_12_7_en( T199 ),
       .io_VwirePorts_0_12_7_out( VwireModule_io_VwirePorts_0_12_7_out ),
       .io_VwirePorts_0_12_6_in( ArrayRowModule_io_V_wire_out_198 ),
       .io_VwirePorts_0_12_6_en( T198 ),
       .io_VwirePorts_0_12_6_out( VwireModule_io_VwirePorts_0_12_6_out ),
       .io_VwirePorts_0_12_5_in( ArrayRowModule_io_V_wire_out_197 ),
       .io_VwirePorts_0_12_5_en( T197 ),
       .io_VwirePorts_0_12_5_out( VwireModule_io_VwirePorts_0_12_5_out ),
       .io_VwirePorts_0_12_4_in( ArrayRowModule_io_V_wire_out_196 ),
       .io_VwirePorts_0_12_4_en( T196 ),
       .io_VwirePorts_0_12_4_out( VwireModule_io_VwirePorts_0_12_4_out ),
       .io_VwirePorts_0_12_3_in( ArrayRowModule_io_V_wire_out_195 ),
       .io_VwirePorts_0_12_3_en( T195 ),
       .io_VwirePorts_0_12_3_out( VwireModule_io_VwirePorts_0_12_3_out ),
       .io_VwirePorts_0_12_2_in( ArrayRowModule_io_V_wire_out_194 ),
       .io_VwirePorts_0_12_2_en( T194 ),
       .io_VwirePorts_0_12_2_out( VwireModule_io_VwirePorts_0_12_2_out ),
       .io_VwirePorts_0_12_1_in( ArrayRowModule_io_V_wire_out_193 ),
       .io_VwirePorts_0_12_1_en( T193 ),
       .io_VwirePorts_0_12_1_out( VwireModule_io_VwirePorts_0_12_1_out ),
       .io_VwirePorts_0_12_0_in( ArrayRowModule_io_V_wire_out_192 ),
       .io_VwirePorts_0_12_0_en( T192 ),
       .io_VwirePorts_0_12_0_out( VwireModule_io_VwirePorts_0_12_0_out ),
       .io_VwirePorts_0_11_15_in( ArrayRowModule_io_V_wire_out_191 ),
       .io_VwirePorts_0_11_15_en( T191 ),
       .io_VwirePorts_0_11_15_out( VwireModule_io_VwirePorts_0_11_15_out ),
       .io_VwirePorts_0_11_14_in( ArrayRowModule_io_V_wire_out_190 ),
       .io_VwirePorts_0_11_14_en( T190 ),
       .io_VwirePorts_0_11_14_out( VwireModule_io_VwirePorts_0_11_14_out ),
       .io_VwirePorts_0_11_13_in( ArrayRowModule_io_V_wire_out_189 ),
       .io_VwirePorts_0_11_13_en( T189 ),
       .io_VwirePorts_0_11_13_out( VwireModule_io_VwirePorts_0_11_13_out ),
       .io_VwirePorts_0_11_12_in( ArrayRowModule_io_V_wire_out_188 ),
       .io_VwirePorts_0_11_12_en( T188 ),
       .io_VwirePorts_0_11_12_out( VwireModule_io_VwirePorts_0_11_12_out ),
       .io_VwirePorts_0_11_11_in( ArrayRowModule_io_V_wire_out_187 ),
       .io_VwirePorts_0_11_11_en( T187 ),
       .io_VwirePorts_0_11_11_out( VwireModule_io_VwirePorts_0_11_11_out ),
       .io_VwirePorts_0_11_10_in( ArrayRowModule_io_V_wire_out_186 ),
       .io_VwirePorts_0_11_10_en( T186 ),
       .io_VwirePorts_0_11_10_out( VwireModule_io_VwirePorts_0_11_10_out ),
       .io_VwirePorts_0_11_9_in( ArrayRowModule_io_V_wire_out_185 ),
       .io_VwirePorts_0_11_9_en( T185 ),
       .io_VwirePorts_0_11_9_out( VwireModule_io_VwirePorts_0_11_9_out ),
       .io_VwirePorts_0_11_8_in( ArrayRowModule_io_V_wire_out_184 ),
       .io_VwirePorts_0_11_8_en( T184 ),
       .io_VwirePorts_0_11_8_out( VwireModule_io_VwirePorts_0_11_8_out ),
       .io_VwirePorts_0_11_7_in( ArrayRowModule_io_V_wire_out_183 ),
       .io_VwirePorts_0_11_7_en( T183 ),
       .io_VwirePorts_0_11_7_out( VwireModule_io_VwirePorts_0_11_7_out ),
       .io_VwirePorts_0_11_6_in( ArrayRowModule_io_V_wire_out_182 ),
       .io_VwirePorts_0_11_6_en( T182 ),
       .io_VwirePorts_0_11_6_out( VwireModule_io_VwirePorts_0_11_6_out ),
       .io_VwirePorts_0_11_5_in( ArrayRowModule_io_V_wire_out_181 ),
       .io_VwirePorts_0_11_5_en( T181 ),
       .io_VwirePorts_0_11_5_out( VwireModule_io_VwirePorts_0_11_5_out ),
       .io_VwirePorts_0_11_4_in( ArrayRowModule_io_V_wire_out_180 ),
       .io_VwirePorts_0_11_4_en( T180 ),
       .io_VwirePorts_0_11_4_out( VwireModule_io_VwirePorts_0_11_4_out ),
       .io_VwirePorts_0_11_3_in( ArrayRowModule_io_V_wire_out_179 ),
       .io_VwirePorts_0_11_3_en( T179 ),
       .io_VwirePorts_0_11_3_out( VwireModule_io_VwirePorts_0_11_3_out ),
       .io_VwirePorts_0_11_2_in( ArrayRowModule_io_V_wire_out_178 ),
       .io_VwirePorts_0_11_2_en( T178 ),
       .io_VwirePorts_0_11_2_out( VwireModule_io_VwirePorts_0_11_2_out ),
       .io_VwirePorts_0_11_1_in( ArrayRowModule_io_V_wire_out_177 ),
       .io_VwirePorts_0_11_1_en( T177 ),
       .io_VwirePorts_0_11_1_out( VwireModule_io_VwirePorts_0_11_1_out ),
       .io_VwirePorts_0_11_0_in( ArrayRowModule_io_V_wire_out_176 ),
       .io_VwirePorts_0_11_0_en( T176 ),
       .io_VwirePorts_0_11_0_out( VwireModule_io_VwirePorts_0_11_0_out ),
       .io_VwirePorts_0_10_15_in( ArrayRowModule_io_V_wire_out_175 ),
       .io_VwirePorts_0_10_15_en( T175 ),
       .io_VwirePorts_0_10_15_out( VwireModule_io_VwirePorts_0_10_15_out ),
       .io_VwirePorts_0_10_14_in( ArrayRowModule_io_V_wire_out_174 ),
       .io_VwirePorts_0_10_14_en( T174 ),
       .io_VwirePorts_0_10_14_out( VwireModule_io_VwirePorts_0_10_14_out ),
       .io_VwirePorts_0_10_13_in( ArrayRowModule_io_V_wire_out_173 ),
       .io_VwirePorts_0_10_13_en( T173 ),
       .io_VwirePorts_0_10_13_out( VwireModule_io_VwirePorts_0_10_13_out ),
       .io_VwirePorts_0_10_12_in( ArrayRowModule_io_V_wire_out_172 ),
       .io_VwirePorts_0_10_12_en( T172 ),
       .io_VwirePorts_0_10_12_out( VwireModule_io_VwirePorts_0_10_12_out ),
       .io_VwirePorts_0_10_11_in( ArrayRowModule_io_V_wire_out_171 ),
       .io_VwirePorts_0_10_11_en( T171 ),
       .io_VwirePorts_0_10_11_out( VwireModule_io_VwirePorts_0_10_11_out ),
       .io_VwirePorts_0_10_10_in( ArrayRowModule_io_V_wire_out_170 ),
       .io_VwirePorts_0_10_10_en( T170 ),
       .io_VwirePorts_0_10_10_out( VwireModule_io_VwirePorts_0_10_10_out ),
       .io_VwirePorts_0_10_9_in( ArrayRowModule_io_V_wire_out_169 ),
       .io_VwirePorts_0_10_9_en( T169 ),
       .io_VwirePorts_0_10_9_out( VwireModule_io_VwirePorts_0_10_9_out ),
       .io_VwirePorts_0_10_8_in( ArrayRowModule_io_V_wire_out_168 ),
       .io_VwirePorts_0_10_8_en( T168 ),
       .io_VwirePorts_0_10_8_out( VwireModule_io_VwirePorts_0_10_8_out ),
       .io_VwirePorts_0_10_7_in( ArrayRowModule_io_V_wire_out_167 ),
       .io_VwirePorts_0_10_7_en( T167 ),
       .io_VwirePorts_0_10_7_out( VwireModule_io_VwirePorts_0_10_7_out ),
       .io_VwirePorts_0_10_6_in( ArrayRowModule_io_V_wire_out_166 ),
       .io_VwirePorts_0_10_6_en( T166 ),
       .io_VwirePorts_0_10_6_out( VwireModule_io_VwirePorts_0_10_6_out ),
       .io_VwirePorts_0_10_5_in( ArrayRowModule_io_V_wire_out_165 ),
       .io_VwirePorts_0_10_5_en( T165 ),
       .io_VwirePorts_0_10_5_out( VwireModule_io_VwirePorts_0_10_5_out ),
       .io_VwirePorts_0_10_4_in( ArrayRowModule_io_V_wire_out_164 ),
       .io_VwirePorts_0_10_4_en( T164 ),
       .io_VwirePorts_0_10_4_out( VwireModule_io_VwirePorts_0_10_4_out ),
       .io_VwirePorts_0_10_3_in( ArrayRowModule_io_V_wire_out_163 ),
       .io_VwirePorts_0_10_3_en( T163 ),
       .io_VwirePorts_0_10_3_out( VwireModule_io_VwirePorts_0_10_3_out ),
       .io_VwirePorts_0_10_2_in( ArrayRowModule_io_V_wire_out_162 ),
       .io_VwirePorts_0_10_2_en( T162 ),
       .io_VwirePorts_0_10_2_out( VwireModule_io_VwirePorts_0_10_2_out ),
       .io_VwirePorts_0_10_1_in( ArrayRowModule_io_V_wire_out_161 ),
       .io_VwirePorts_0_10_1_en( T161 ),
       .io_VwirePorts_0_10_1_out( VwireModule_io_VwirePorts_0_10_1_out ),
       .io_VwirePorts_0_10_0_in( ArrayRowModule_io_V_wire_out_160 ),
       .io_VwirePorts_0_10_0_en( T160 ),
       .io_VwirePorts_0_10_0_out( VwireModule_io_VwirePorts_0_10_0_out ),
       .io_VwirePorts_0_9_15_in( ArrayRowModule_io_V_wire_out_159 ),
       .io_VwirePorts_0_9_15_en( T159 ),
       .io_VwirePorts_0_9_15_out( VwireModule_io_VwirePorts_0_9_15_out ),
       .io_VwirePorts_0_9_14_in( ArrayRowModule_io_V_wire_out_158 ),
       .io_VwirePorts_0_9_14_en( T158 ),
       .io_VwirePorts_0_9_14_out( VwireModule_io_VwirePorts_0_9_14_out ),
       .io_VwirePorts_0_9_13_in( ArrayRowModule_io_V_wire_out_157 ),
       .io_VwirePorts_0_9_13_en( T157 ),
       .io_VwirePorts_0_9_13_out( VwireModule_io_VwirePorts_0_9_13_out ),
       .io_VwirePorts_0_9_12_in( ArrayRowModule_io_V_wire_out_156 ),
       .io_VwirePorts_0_9_12_en( T156 ),
       .io_VwirePorts_0_9_12_out( VwireModule_io_VwirePorts_0_9_12_out ),
       .io_VwirePorts_0_9_11_in( ArrayRowModule_io_V_wire_out_155 ),
       .io_VwirePorts_0_9_11_en( T155 ),
       .io_VwirePorts_0_9_11_out( VwireModule_io_VwirePorts_0_9_11_out ),
       .io_VwirePorts_0_9_10_in( ArrayRowModule_io_V_wire_out_154 ),
       .io_VwirePorts_0_9_10_en( T154 ),
       .io_VwirePorts_0_9_10_out( VwireModule_io_VwirePorts_0_9_10_out ),
       .io_VwirePorts_0_9_9_in( ArrayRowModule_io_V_wire_out_153 ),
       .io_VwirePorts_0_9_9_en( T153 ),
       .io_VwirePorts_0_9_9_out( VwireModule_io_VwirePorts_0_9_9_out ),
       .io_VwirePorts_0_9_8_in( ArrayRowModule_io_V_wire_out_152 ),
       .io_VwirePorts_0_9_8_en( T152 ),
       .io_VwirePorts_0_9_8_out( VwireModule_io_VwirePorts_0_9_8_out ),
       .io_VwirePorts_0_9_7_in( ArrayRowModule_io_V_wire_out_151 ),
       .io_VwirePorts_0_9_7_en( T151 ),
       .io_VwirePorts_0_9_7_out( VwireModule_io_VwirePorts_0_9_7_out ),
       .io_VwirePorts_0_9_6_in( ArrayRowModule_io_V_wire_out_150 ),
       .io_VwirePorts_0_9_6_en( T150 ),
       .io_VwirePorts_0_9_6_out( VwireModule_io_VwirePorts_0_9_6_out ),
       .io_VwirePorts_0_9_5_in( ArrayRowModule_io_V_wire_out_149 ),
       .io_VwirePorts_0_9_5_en( T149 ),
       .io_VwirePorts_0_9_5_out( VwireModule_io_VwirePorts_0_9_5_out ),
       .io_VwirePorts_0_9_4_in( ArrayRowModule_io_V_wire_out_148 ),
       .io_VwirePorts_0_9_4_en( T148 ),
       .io_VwirePorts_0_9_4_out( VwireModule_io_VwirePorts_0_9_4_out ),
       .io_VwirePorts_0_9_3_in( ArrayRowModule_io_V_wire_out_147 ),
       .io_VwirePorts_0_9_3_en( T147 ),
       .io_VwirePorts_0_9_3_out( VwireModule_io_VwirePorts_0_9_3_out ),
       .io_VwirePorts_0_9_2_in( ArrayRowModule_io_V_wire_out_146 ),
       .io_VwirePorts_0_9_2_en( T146 ),
       .io_VwirePorts_0_9_2_out( VwireModule_io_VwirePorts_0_9_2_out ),
       .io_VwirePorts_0_9_1_in( ArrayRowModule_io_V_wire_out_145 ),
       .io_VwirePorts_0_9_1_en( T145 ),
       .io_VwirePorts_0_9_1_out( VwireModule_io_VwirePorts_0_9_1_out ),
       .io_VwirePorts_0_9_0_in( ArrayRowModule_io_V_wire_out_144 ),
       .io_VwirePorts_0_9_0_en( T144 ),
       .io_VwirePorts_0_9_0_out( VwireModule_io_VwirePorts_0_9_0_out ),
       .io_VwirePorts_0_8_15_in( ArrayRowModule_io_V_wire_out_143 ),
       .io_VwirePorts_0_8_15_en( T143 ),
       .io_VwirePorts_0_8_15_out( VwireModule_io_VwirePorts_0_8_15_out ),
       .io_VwirePorts_0_8_14_in( ArrayRowModule_io_V_wire_out_142 ),
       .io_VwirePorts_0_8_14_en( T142 ),
       .io_VwirePorts_0_8_14_out( VwireModule_io_VwirePorts_0_8_14_out ),
       .io_VwirePorts_0_8_13_in( ArrayRowModule_io_V_wire_out_141 ),
       .io_VwirePorts_0_8_13_en( T141 ),
       .io_VwirePorts_0_8_13_out( VwireModule_io_VwirePorts_0_8_13_out ),
       .io_VwirePorts_0_8_12_in( ArrayRowModule_io_V_wire_out_140 ),
       .io_VwirePorts_0_8_12_en( T140 ),
       .io_VwirePorts_0_8_12_out( VwireModule_io_VwirePorts_0_8_12_out ),
       .io_VwirePorts_0_8_11_in( ArrayRowModule_io_V_wire_out_139 ),
       .io_VwirePorts_0_8_11_en( T139 ),
       .io_VwirePorts_0_8_11_out( VwireModule_io_VwirePorts_0_8_11_out ),
       .io_VwirePorts_0_8_10_in( ArrayRowModule_io_V_wire_out_138 ),
       .io_VwirePorts_0_8_10_en( T138 ),
       .io_VwirePorts_0_8_10_out( VwireModule_io_VwirePorts_0_8_10_out ),
       .io_VwirePorts_0_8_9_in( ArrayRowModule_io_V_wire_out_137 ),
       .io_VwirePorts_0_8_9_en( T137 ),
       .io_VwirePorts_0_8_9_out( VwireModule_io_VwirePorts_0_8_9_out ),
       .io_VwirePorts_0_8_8_in( ArrayRowModule_io_V_wire_out_136 ),
       .io_VwirePorts_0_8_8_en( T136 ),
       .io_VwirePorts_0_8_8_out( VwireModule_io_VwirePorts_0_8_8_out ),
       .io_VwirePorts_0_8_7_in( ArrayRowModule_io_V_wire_out_135 ),
       .io_VwirePorts_0_8_7_en( T135 ),
       .io_VwirePorts_0_8_7_out( VwireModule_io_VwirePorts_0_8_7_out ),
       .io_VwirePorts_0_8_6_in( ArrayRowModule_io_V_wire_out_134 ),
       .io_VwirePorts_0_8_6_en( T134 ),
       .io_VwirePorts_0_8_6_out( VwireModule_io_VwirePorts_0_8_6_out ),
       .io_VwirePorts_0_8_5_in( ArrayRowModule_io_V_wire_out_133 ),
       .io_VwirePorts_0_8_5_en( T133 ),
       .io_VwirePorts_0_8_5_out( VwireModule_io_VwirePorts_0_8_5_out ),
       .io_VwirePorts_0_8_4_in( ArrayRowModule_io_V_wire_out_132 ),
       .io_VwirePorts_0_8_4_en( T132 ),
       .io_VwirePorts_0_8_4_out( VwireModule_io_VwirePorts_0_8_4_out ),
       .io_VwirePorts_0_8_3_in( ArrayRowModule_io_V_wire_out_131 ),
       .io_VwirePorts_0_8_3_en( T131 ),
       .io_VwirePorts_0_8_3_out( VwireModule_io_VwirePorts_0_8_3_out ),
       .io_VwirePorts_0_8_2_in( ArrayRowModule_io_V_wire_out_130 ),
       .io_VwirePorts_0_8_2_en( T130 ),
       .io_VwirePorts_0_8_2_out( VwireModule_io_VwirePorts_0_8_2_out ),
       .io_VwirePorts_0_8_1_in( ArrayRowModule_io_V_wire_out_129 ),
       .io_VwirePorts_0_8_1_en( T129 ),
       .io_VwirePorts_0_8_1_out( VwireModule_io_VwirePorts_0_8_1_out ),
       .io_VwirePorts_0_8_0_in( ArrayRowModule_io_V_wire_out_128 ),
       .io_VwirePorts_0_8_0_en( T128 ),
       .io_VwirePorts_0_8_0_out( VwireModule_io_VwirePorts_0_8_0_out ),
       .io_VwirePorts_0_7_15_in( ArrayRowModule_io_V_wire_out_127 ),
       .io_VwirePorts_0_7_15_en( T127 ),
       .io_VwirePorts_0_7_15_out( VwireModule_io_VwirePorts_0_7_15_out ),
       .io_VwirePorts_0_7_14_in( ArrayRowModule_io_V_wire_out_126 ),
       .io_VwirePorts_0_7_14_en( T126 ),
       .io_VwirePorts_0_7_14_out( VwireModule_io_VwirePorts_0_7_14_out ),
       .io_VwirePorts_0_7_13_in( ArrayRowModule_io_V_wire_out_125 ),
       .io_VwirePorts_0_7_13_en( T125 ),
       .io_VwirePorts_0_7_13_out( VwireModule_io_VwirePorts_0_7_13_out ),
       .io_VwirePorts_0_7_12_in( ArrayRowModule_io_V_wire_out_124 ),
       .io_VwirePorts_0_7_12_en( T124 ),
       .io_VwirePorts_0_7_12_out( VwireModule_io_VwirePorts_0_7_12_out ),
       .io_VwirePorts_0_7_11_in( ArrayRowModule_io_V_wire_out_123 ),
       .io_VwirePorts_0_7_11_en( T123 ),
       .io_VwirePorts_0_7_11_out( VwireModule_io_VwirePorts_0_7_11_out ),
       .io_VwirePorts_0_7_10_in( ArrayRowModule_io_V_wire_out_122 ),
       .io_VwirePorts_0_7_10_en( T122 ),
       .io_VwirePorts_0_7_10_out( VwireModule_io_VwirePorts_0_7_10_out ),
       .io_VwirePorts_0_7_9_in( ArrayRowModule_io_V_wire_out_121 ),
       .io_VwirePorts_0_7_9_en( T121 ),
       .io_VwirePorts_0_7_9_out( VwireModule_io_VwirePorts_0_7_9_out ),
       .io_VwirePorts_0_7_8_in( ArrayRowModule_io_V_wire_out_120 ),
       .io_VwirePorts_0_7_8_en( T120 ),
       .io_VwirePorts_0_7_8_out( VwireModule_io_VwirePorts_0_7_8_out ),
       .io_VwirePorts_0_7_7_in( ArrayRowModule_io_V_wire_out_119 ),
       .io_VwirePorts_0_7_7_en( T119 ),
       .io_VwirePorts_0_7_7_out( VwireModule_io_VwirePorts_0_7_7_out ),
       .io_VwirePorts_0_7_6_in( ArrayRowModule_io_V_wire_out_118 ),
       .io_VwirePorts_0_7_6_en( T118 ),
       .io_VwirePorts_0_7_6_out( VwireModule_io_VwirePorts_0_7_6_out ),
       .io_VwirePorts_0_7_5_in( ArrayRowModule_io_V_wire_out_117 ),
       .io_VwirePorts_0_7_5_en( T117 ),
       .io_VwirePorts_0_7_5_out( VwireModule_io_VwirePorts_0_7_5_out ),
       .io_VwirePorts_0_7_4_in( ArrayRowModule_io_V_wire_out_116 ),
       .io_VwirePorts_0_7_4_en( T116 ),
       .io_VwirePorts_0_7_4_out( VwireModule_io_VwirePorts_0_7_4_out ),
       .io_VwirePorts_0_7_3_in( ArrayRowModule_io_V_wire_out_115 ),
       .io_VwirePorts_0_7_3_en( T115 ),
       .io_VwirePorts_0_7_3_out( VwireModule_io_VwirePorts_0_7_3_out ),
       .io_VwirePorts_0_7_2_in( ArrayRowModule_io_V_wire_out_114 ),
       .io_VwirePorts_0_7_2_en( T114 ),
       .io_VwirePorts_0_7_2_out( VwireModule_io_VwirePorts_0_7_2_out ),
       .io_VwirePorts_0_7_1_in( ArrayRowModule_io_V_wire_out_113 ),
       .io_VwirePorts_0_7_1_en( T113 ),
       .io_VwirePorts_0_7_1_out( VwireModule_io_VwirePorts_0_7_1_out ),
       .io_VwirePorts_0_7_0_in( ArrayRowModule_io_V_wire_out_112 ),
       .io_VwirePorts_0_7_0_en( T112 ),
       .io_VwirePorts_0_7_0_out( VwireModule_io_VwirePorts_0_7_0_out ),
       .io_VwirePorts_0_6_15_in( ArrayRowModule_io_V_wire_out_111 ),
       .io_VwirePorts_0_6_15_en( T111 ),
       .io_VwirePorts_0_6_15_out( VwireModule_io_VwirePorts_0_6_15_out ),
       .io_VwirePorts_0_6_14_in( ArrayRowModule_io_V_wire_out_110 ),
       .io_VwirePorts_0_6_14_en( T110 ),
       .io_VwirePorts_0_6_14_out( VwireModule_io_VwirePorts_0_6_14_out ),
       .io_VwirePorts_0_6_13_in( ArrayRowModule_io_V_wire_out_109 ),
       .io_VwirePorts_0_6_13_en( T109 ),
       .io_VwirePorts_0_6_13_out( VwireModule_io_VwirePorts_0_6_13_out ),
       .io_VwirePorts_0_6_12_in( ArrayRowModule_io_V_wire_out_108 ),
       .io_VwirePorts_0_6_12_en( T108 ),
       .io_VwirePorts_0_6_12_out( VwireModule_io_VwirePorts_0_6_12_out ),
       .io_VwirePorts_0_6_11_in( ArrayRowModule_io_V_wire_out_107 ),
       .io_VwirePorts_0_6_11_en( T107 ),
       .io_VwirePorts_0_6_11_out( VwireModule_io_VwirePorts_0_6_11_out ),
       .io_VwirePorts_0_6_10_in( ArrayRowModule_io_V_wire_out_106 ),
       .io_VwirePorts_0_6_10_en( T106 ),
       .io_VwirePorts_0_6_10_out( VwireModule_io_VwirePorts_0_6_10_out ),
       .io_VwirePorts_0_6_9_in( ArrayRowModule_io_V_wire_out_105 ),
       .io_VwirePorts_0_6_9_en( T105 ),
       .io_VwirePorts_0_6_9_out( VwireModule_io_VwirePorts_0_6_9_out ),
       .io_VwirePorts_0_6_8_in( ArrayRowModule_io_V_wire_out_104 ),
       .io_VwirePorts_0_6_8_en( T104 ),
       .io_VwirePorts_0_6_8_out( VwireModule_io_VwirePorts_0_6_8_out ),
       .io_VwirePorts_0_6_7_in( ArrayRowModule_io_V_wire_out_103 ),
       .io_VwirePorts_0_6_7_en( T103 ),
       .io_VwirePorts_0_6_7_out( VwireModule_io_VwirePorts_0_6_7_out ),
       .io_VwirePorts_0_6_6_in( ArrayRowModule_io_V_wire_out_102 ),
       .io_VwirePorts_0_6_6_en( T102 ),
       .io_VwirePorts_0_6_6_out( VwireModule_io_VwirePorts_0_6_6_out ),
       .io_VwirePorts_0_6_5_in( ArrayRowModule_io_V_wire_out_101 ),
       .io_VwirePorts_0_6_5_en( T101 ),
       .io_VwirePorts_0_6_5_out( VwireModule_io_VwirePorts_0_6_5_out ),
       .io_VwirePorts_0_6_4_in( ArrayRowModule_io_V_wire_out_100 ),
       .io_VwirePorts_0_6_4_en( T100 ),
       .io_VwirePorts_0_6_4_out( VwireModule_io_VwirePorts_0_6_4_out ),
       .io_VwirePorts_0_6_3_in( ArrayRowModule_io_V_wire_out_99 ),
       .io_VwirePorts_0_6_3_en( T99 ),
       .io_VwirePorts_0_6_3_out( VwireModule_io_VwirePorts_0_6_3_out ),
       .io_VwirePorts_0_6_2_in( ArrayRowModule_io_V_wire_out_98 ),
       .io_VwirePorts_0_6_2_en( T98 ),
       .io_VwirePorts_0_6_2_out( VwireModule_io_VwirePorts_0_6_2_out ),
       .io_VwirePorts_0_6_1_in( ArrayRowModule_io_V_wire_out_97 ),
       .io_VwirePorts_0_6_1_en( T97 ),
       .io_VwirePorts_0_6_1_out( VwireModule_io_VwirePorts_0_6_1_out ),
       .io_VwirePorts_0_6_0_in( ArrayRowModule_io_V_wire_out_96 ),
       .io_VwirePorts_0_6_0_en( T96 ),
       .io_VwirePorts_0_6_0_out( VwireModule_io_VwirePorts_0_6_0_out ),
       .io_VwirePorts_0_5_15_in( ArrayRowModule_io_V_wire_out_95 ),
       .io_VwirePorts_0_5_15_en( T95 ),
       .io_VwirePorts_0_5_15_out( VwireModule_io_VwirePorts_0_5_15_out ),
       .io_VwirePorts_0_5_14_in( ArrayRowModule_io_V_wire_out_94 ),
       .io_VwirePorts_0_5_14_en( T94 ),
       .io_VwirePorts_0_5_14_out( VwireModule_io_VwirePorts_0_5_14_out ),
       .io_VwirePorts_0_5_13_in( ArrayRowModule_io_V_wire_out_93 ),
       .io_VwirePorts_0_5_13_en( T93 ),
       .io_VwirePorts_0_5_13_out( VwireModule_io_VwirePorts_0_5_13_out ),
       .io_VwirePorts_0_5_12_in( ArrayRowModule_io_V_wire_out_92 ),
       .io_VwirePorts_0_5_12_en( T92 ),
       .io_VwirePorts_0_5_12_out( VwireModule_io_VwirePorts_0_5_12_out ),
       .io_VwirePorts_0_5_11_in( ArrayRowModule_io_V_wire_out_91 ),
       .io_VwirePorts_0_5_11_en( T91 ),
       .io_VwirePorts_0_5_11_out( VwireModule_io_VwirePorts_0_5_11_out ),
       .io_VwirePorts_0_5_10_in( ArrayRowModule_io_V_wire_out_90 ),
       .io_VwirePorts_0_5_10_en( T90 ),
       .io_VwirePorts_0_5_10_out( VwireModule_io_VwirePorts_0_5_10_out ),
       .io_VwirePorts_0_5_9_in( ArrayRowModule_io_V_wire_out_89 ),
       .io_VwirePorts_0_5_9_en( T89 ),
       .io_VwirePorts_0_5_9_out( VwireModule_io_VwirePorts_0_5_9_out ),
       .io_VwirePorts_0_5_8_in( ArrayRowModule_io_V_wire_out_88 ),
       .io_VwirePorts_0_5_8_en( T88 ),
       .io_VwirePorts_0_5_8_out( VwireModule_io_VwirePorts_0_5_8_out ),
       .io_VwirePorts_0_5_7_in( ArrayRowModule_io_V_wire_out_87 ),
       .io_VwirePorts_0_5_7_en( T87 ),
       .io_VwirePorts_0_5_7_out( VwireModule_io_VwirePorts_0_5_7_out ),
       .io_VwirePorts_0_5_6_in( ArrayRowModule_io_V_wire_out_86 ),
       .io_VwirePorts_0_5_6_en( T86 ),
       .io_VwirePorts_0_5_6_out( VwireModule_io_VwirePorts_0_5_6_out ),
       .io_VwirePorts_0_5_5_in( ArrayRowModule_io_V_wire_out_85 ),
       .io_VwirePorts_0_5_5_en( T85 ),
       .io_VwirePorts_0_5_5_out( VwireModule_io_VwirePorts_0_5_5_out ),
       .io_VwirePorts_0_5_4_in( ArrayRowModule_io_V_wire_out_84 ),
       .io_VwirePorts_0_5_4_en( T84 ),
       .io_VwirePorts_0_5_4_out( VwireModule_io_VwirePorts_0_5_4_out ),
       .io_VwirePorts_0_5_3_in( ArrayRowModule_io_V_wire_out_83 ),
       .io_VwirePorts_0_5_3_en( T83 ),
       .io_VwirePorts_0_5_3_out( VwireModule_io_VwirePorts_0_5_3_out ),
       .io_VwirePorts_0_5_2_in( ArrayRowModule_io_V_wire_out_82 ),
       .io_VwirePorts_0_5_2_en( T82 ),
       .io_VwirePorts_0_5_2_out( VwireModule_io_VwirePorts_0_5_2_out ),
       .io_VwirePorts_0_5_1_in( ArrayRowModule_io_V_wire_out_81 ),
       .io_VwirePorts_0_5_1_en( T81 ),
       .io_VwirePorts_0_5_1_out( VwireModule_io_VwirePorts_0_5_1_out ),
       .io_VwirePorts_0_5_0_in( ArrayRowModule_io_V_wire_out_80 ),
       .io_VwirePorts_0_5_0_en( T80 ),
       .io_VwirePorts_0_5_0_out( VwireModule_io_VwirePorts_0_5_0_out ),
       .io_VwirePorts_0_4_15_in( ArrayRowModule_io_V_wire_out_79 ),
       .io_VwirePorts_0_4_15_en( T79 ),
       .io_VwirePorts_0_4_15_out( VwireModule_io_VwirePorts_0_4_15_out ),
       .io_VwirePorts_0_4_14_in( ArrayRowModule_io_V_wire_out_78 ),
       .io_VwirePorts_0_4_14_en( T78 ),
       .io_VwirePorts_0_4_14_out( VwireModule_io_VwirePorts_0_4_14_out ),
       .io_VwirePorts_0_4_13_in( ArrayRowModule_io_V_wire_out_77 ),
       .io_VwirePorts_0_4_13_en( T77 ),
       .io_VwirePorts_0_4_13_out( VwireModule_io_VwirePorts_0_4_13_out ),
       .io_VwirePorts_0_4_12_in( ArrayRowModule_io_V_wire_out_76 ),
       .io_VwirePorts_0_4_12_en( T76 ),
       .io_VwirePorts_0_4_12_out( VwireModule_io_VwirePorts_0_4_12_out ),
       .io_VwirePorts_0_4_11_in( ArrayRowModule_io_V_wire_out_75 ),
       .io_VwirePorts_0_4_11_en( T75 ),
       .io_VwirePorts_0_4_11_out( VwireModule_io_VwirePorts_0_4_11_out ),
       .io_VwirePorts_0_4_10_in( ArrayRowModule_io_V_wire_out_74 ),
       .io_VwirePorts_0_4_10_en( T74 ),
       .io_VwirePorts_0_4_10_out( VwireModule_io_VwirePorts_0_4_10_out ),
       .io_VwirePorts_0_4_9_in( ArrayRowModule_io_V_wire_out_73 ),
       .io_VwirePorts_0_4_9_en( T73 ),
       .io_VwirePorts_0_4_9_out( VwireModule_io_VwirePorts_0_4_9_out ),
       .io_VwirePorts_0_4_8_in( ArrayRowModule_io_V_wire_out_72 ),
       .io_VwirePorts_0_4_8_en( T72 ),
       .io_VwirePorts_0_4_8_out( VwireModule_io_VwirePorts_0_4_8_out ),
       .io_VwirePorts_0_4_7_in( ArrayRowModule_io_V_wire_out_71 ),
       .io_VwirePorts_0_4_7_en( T71 ),
       .io_VwirePorts_0_4_7_out( VwireModule_io_VwirePorts_0_4_7_out ),
       .io_VwirePorts_0_4_6_in( ArrayRowModule_io_V_wire_out_70 ),
       .io_VwirePorts_0_4_6_en( T70 ),
       .io_VwirePorts_0_4_6_out( VwireModule_io_VwirePorts_0_4_6_out ),
       .io_VwirePorts_0_4_5_in( ArrayRowModule_io_V_wire_out_69 ),
       .io_VwirePorts_0_4_5_en( T69 ),
       .io_VwirePorts_0_4_5_out( VwireModule_io_VwirePorts_0_4_5_out ),
       .io_VwirePorts_0_4_4_in( ArrayRowModule_io_V_wire_out_68 ),
       .io_VwirePorts_0_4_4_en( T68 ),
       .io_VwirePorts_0_4_4_out( VwireModule_io_VwirePorts_0_4_4_out ),
       .io_VwirePorts_0_4_3_in( ArrayRowModule_io_V_wire_out_67 ),
       .io_VwirePorts_0_4_3_en( T67 ),
       .io_VwirePorts_0_4_3_out( VwireModule_io_VwirePorts_0_4_3_out ),
       .io_VwirePorts_0_4_2_in( ArrayRowModule_io_V_wire_out_66 ),
       .io_VwirePorts_0_4_2_en( T66 ),
       .io_VwirePorts_0_4_2_out( VwireModule_io_VwirePorts_0_4_2_out ),
       .io_VwirePorts_0_4_1_in( ArrayRowModule_io_V_wire_out_65 ),
       .io_VwirePorts_0_4_1_en( T65 ),
       .io_VwirePorts_0_4_1_out( VwireModule_io_VwirePorts_0_4_1_out ),
       .io_VwirePorts_0_4_0_in( ArrayRowModule_io_V_wire_out_64 ),
       .io_VwirePorts_0_4_0_en( T64 ),
       .io_VwirePorts_0_4_0_out( VwireModule_io_VwirePorts_0_4_0_out ),
       .io_VwirePorts_0_3_15_in( ArrayRowModule_io_V_wire_out_63 ),
       .io_VwirePorts_0_3_15_en( T63 ),
       .io_VwirePorts_0_3_15_out( VwireModule_io_VwirePorts_0_3_15_out ),
       .io_VwirePorts_0_3_14_in( ArrayRowModule_io_V_wire_out_62 ),
       .io_VwirePorts_0_3_14_en( T62 ),
       .io_VwirePorts_0_3_14_out( VwireModule_io_VwirePorts_0_3_14_out ),
       .io_VwirePorts_0_3_13_in( ArrayRowModule_io_V_wire_out_61 ),
       .io_VwirePorts_0_3_13_en( T61 ),
       .io_VwirePorts_0_3_13_out( VwireModule_io_VwirePorts_0_3_13_out ),
       .io_VwirePorts_0_3_12_in( ArrayRowModule_io_V_wire_out_60 ),
       .io_VwirePorts_0_3_12_en( T60 ),
       .io_VwirePorts_0_3_12_out( VwireModule_io_VwirePorts_0_3_12_out ),
       .io_VwirePorts_0_3_11_in( ArrayRowModule_io_V_wire_out_59 ),
       .io_VwirePorts_0_3_11_en( T59 ),
       .io_VwirePorts_0_3_11_out( VwireModule_io_VwirePorts_0_3_11_out ),
       .io_VwirePorts_0_3_10_in( ArrayRowModule_io_V_wire_out_58 ),
       .io_VwirePorts_0_3_10_en( T58 ),
       .io_VwirePorts_0_3_10_out( VwireModule_io_VwirePorts_0_3_10_out ),
       .io_VwirePorts_0_3_9_in( ArrayRowModule_io_V_wire_out_57 ),
       .io_VwirePorts_0_3_9_en( T57 ),
       .io_VwirePorts_0_3_9_out( VwireModule_io_VwirePorts_0_3_9_out ),
       .io_VwirePorts_0_3_8_in( ArrayRowModule_io_V_wire_out_56 ),
       .io_VwirePorts_0_3_8_en( T56 ),
       .io_VwirePorts_0_3_8_out( VwireModule_io_VwirePorts_0_3_8_out ),
       .io_VwirePorts_0_3_7_in( ArrayRowModule_io_V_wire_out_55 ),
       .io_VwirePorts_0_3_7_en( T55 ),
       .io_VwirePorts_0_3_7_out( VwireModule_io_VwirePorts_0_3_7_out ),
       .io_VwirePorts_0_3_6_in( ArrayRowModule_io_V_wire_out_54 ),
       .io_VwirePorts_0_3_6_en( T54 ),
       .io_VwirePorts_0_3_6_out( VwireModule_io_VwirePorts_0_3_6_out ),
       .io_VwirePorts_0_3_5_in( ArrayRowModule_io_V_wire_out_53 ),
       .io_VwirePorts_0_3_5_en( T53 ),
       .io_VwirePorts_0_3_5_out( VwireModule_io_VwirePorts_0_3_5_out ),
       .io_VwirePorts_0_3_4_in( ArrayRowModule_io_V_wire_out_52 ),
       .io_VwirePorts_0_3_4_en( T52 ),
       .io_VwirePorts_0_3_4_out( VwireModule_io_VwirePorts_0_3_4_out ),
       .io_VwirePorts_0_3_3_in( ArrayRowModule_io_V_wire_out_51 ),
       .io_VwirePorts_0_3_3_en( T51 ),
       .io_VwirePorts_0_3_3_out( VwireModule_io_VwirePorts_0_3_3_out ),
       .io_VwirePorts_0_3_2_in( ArrayRowModule_io_V_wire_out_50 ),
       .io_VwirePorts_0_3_2_en( T50 ),
       .io_VwirePorts_0_3_2_out( VwireModule_io_VwirePorts_0_3_2_out ),
       .io_VwirePorts_0_3_1_in( ArrayRowModule_io_V_wire_out_49 ),
       .io_VwirePorts_0_3_1_en( T49 ),
       .io_VwirePorts_0_3_1_out( VwireModule_io_VwirePorts_0_3_1_out ),
       .io_VwirePorts_0_3_0_in( ArrayRowModule_io_V_wire_out_48 ),
       .io_VwirePorts_0_3_0_en( T48 ),
       .io_VwirePorts_0_3_0_out( VwireModule_io_VwirePorts_0_3_0_out ),
       .io_VwirePorts_0_2_15_in( ArrayRowModule_io_V_wire_out_47 ),
       .io_VwirePorts_0_2_15_en( T47 ),
       .io_VwirePorts_0_2_15_out( VwireModule_io_VwirePorts_0_2_15_out ),
       .io_VwirePorts_0_2_14_in( ArrayRowModule_io_V_wire_out_46 ),
       .io_VwirePorts_0_2_14_en( T46 ),
       .io_VwirePorts_0_2_14_out( VwireModule_io_VwirePorts_0_2_14_out ),
       .io_VwirePorts_0_2_13_in( ArrayRowModule_io_V_wire_out_45 ),
       .io_VwirePorts_0_2_13_en( T45 ),
       .io_VwirePorts_0_2_13_out( VwireModule_io_VwirePorts_0_2_13_out ),
       .io_VwirePorts_0_2_12_in( ArrayRowModule_io_V_wire_out_44 ),
       .io_VwirePorts_0_2_12_en( T44 ),
       .io_VwirePorts_0_2_12_out( VwireModule_io_VwirePorts_0_2_12_out ),
       .io_VwirePorts_0_2_11_in( ArrayRowModule_io_V_wire_out_43 ),
       .io_VwirePorts_0_2_11_en( T43 ),
       .io_VwirePorts_0_2_11_out( VwireModule_io_VwirePorts_0_2_11_out ),
       .io_VwirePorts_0_2_10_in( ArrayRowModule_io_V_wire_out_42 ),
       .io_VwirePorts_0_2_10_en( T42 ),
       .io_VwirePorts_0_2_10_out( VwireModule_io_VwirePorts_0_2_10_out ),
       .io_VwirePorts_0_2_9_in( ArrayRowModule_io_V_wire_out_41 ),
       .io_VwirePorts_0_2_9_en( T41 ),
       .io_VwirePorts_0_2_9_out( VwireModule_io_VwirePorts_0_2_9_out ),
       .io_VwirePorts_0_2_8_in( ArrayRowModule_io_V_wire_out_40 ),
       .io_VwirePorts_0_2_8_en( T40 ),
       .io_VwirePorts_0_2_8_out( VwireModule_io_VwirePorts_0_2_8_out ),
       .io_VwirePorts_0_2_7_in( ArrayRowModule_io_V_wire_out_39 ),
       .io_VwirePorts_0_2_7_en( T39 ),
       .io_VwirePorts_0_2_7_out( VwireModule_io_VwirePorts_0_2_7_out ),
       .io_VwirePorts_0_2_6_in( ArrayRowModule_io_V_wire_out_38 ),
       .io_VwirePorts_0_2_6_en( T38 ),
       .io_VwirePorts_0_2_6_out( VwireModule_io_VwirePorts_0_2_6_out ),
       .io_VwirePorts_0_2_5_in( ArrayRowModule_io_V_wire_out_37 ),
       .io_VwirePorts_0_2_5_en( T37 ),
       .io_VwirePorts_0_2_5_out( VwireModule_io_VwirePorts_0_2_5_out ),
       .io_VwirePorts_0_2_4_in( ArrayRowModule_io_V_wire_out_36 ),
       .io_VwirePorts_0_2_4_en( T36 ),
       .io_VwirePorts_0_2_4_out( VwireModule_io_VwirePorts_0_2_4_out ),
       .io_VwirePorts_0_2_3_in( ArrayRowModule_io_V_wire_out_35 ),
       .io_VwirePorts_0_2_3_en( T35 ),
       .io_VwirePorts_0_2_3_out( VwireModule_io_VwirePorts_0_2_3_out ),
       .io_VwirePorts_0_2_2_in( ArrayRowModule_io_V_wire_out_34 ),
       .io_VwirePorts_0_2_2_en( T34 ),
       .io_VwirePorts_0_2_2_out( VwireModule_io_VwirePorts_0_2_2_out ),
       .io_VwirePorts_0_2_1_in( ArrayRowModule_io_V_wire_out_33 ),
       .io_VwirePorts_0_2_1_en( T33 ),
       .io_VwirePorts_0_2_1_out( VwireModule_io_VwirePorts_0_2_1_out ),
       .io_VwirePorts_0_2_0_in( ArrayRowModule_io_V_wire_out_32 ),
       .io_VwirePorts_0_2_0_en( T32 ),
       .io_VwirePorts_0_2_0_out( VwireModule_io_VwirePorts_0_2_0_out ),
       .io_VwirePorts_0_1_15_in( ArrayRowModule_io_V_wire_out_31 ),
       .io_VwirePorts_0_1_15_en( T31 ),
       .io_VwirePorts_0_1_15_out( VwireModule_io_VwirePorts_0_1_15_out ),
       .io_VwirePorts_0_1_14_in( ArrayRowModule_io_V_wire_out_30 ),
       .io_VwirePorts_0_1_14_en( T30 ),
       .io_VwirePorts_0_1_14_out( VwireModule_io_VwirePorts_0_1_14_out ),
       .io_VwirePorts_0_1_13_in( ArrayRowModule_io_V_wire_out_29 ),
       .io_VwirePorts_0_1_13_en( T29 ),
       .io_VwirePorts_0_1_13_out( VwireModule_io_VwirePorts_0_1_13_out ),
       .io_VwirePorts_0_1_12_in( ArrayRowModule_io_V_wire_out_28 ),
       .io_VwirePorts_0_1_12_en( T28 ),
       .io_VwirePorts_0_1_12_out( VwireModule_io_VwirePorts_0_1_12_out ),
       .io_VwirePorts_0_1_11_in( ArrayRowModule_io_V_wire_out_27 ),
       .io_VwirePorts_0_1_11_en( T27 ),
       .io_VwirePorts_0_1_11_out( VwireModule_io_VwirePorts_0_1_11_out ),
       .io_VwirePorts_0_1_10_in( ArrayRowModule_io_V_wire_out_26 ),
       .io_VwirePorts_0_1_10_en( T26 ),
       .io_VwirePorts_0_1_10_out( VwireModule_io_VwirePorts_0_1_10_out ),
       .io_VwirePorts_0_1_9_in( ArrayRowModule_io_V_wire_out_25 ),
       .io_VwirePorts_0_1_9_en( T25 ),
       .io_VwirePorts_0_1_9_out( VwireModule_io_VwirePorts_0_1_9_out ),
       .io_VwirePorts_0_1_8_in( ArrayRowModule_io_V_wire_out_24 ),
       .io_VwirePorts_0_1_8_en( T24 ),
       .io_VwirePorts_0_1_8_out( VwireModule_io_VwirePorts_0_1_8_out ),
       .io_VwirePorts_0_1_7_in( ArrayRowModule_io_V_wire_out_23 ),
       .io_VwirePorts_0_1_7_en( T23 ),
       .io_VwirePorts_0_1_7_out( VwireModule_io_VwirePorts_0_1_7_out ),
       .io_VwirePorts_0_1_6_in( ArrayRowModule_io_V_wire_out_22 ),
       .io_VwirePorts_0_1_6_en( T22 ),
       .io_VwirePorts_0_1_6_out( VwireModule_io_VwirePorts_0_1_6_out ),
       .io_VwirePorts_0_1_5_in( ArrayRowModule_io_V_wire_out_21 ),
       .io_VwirePorts_0_1_5_en( T21 ),
       .io_VwirePorts_0_1_5_out( VwireModule_io_VwirePorts_0_1_5_out ),
       .io_VwirePorts_0_1_4_in( ArrayRowModule_io_V_wire_out_20 ),
       .io_VwirePorts_0_1_4_en( T20 ),
       .io_VwirePorts_0_1_4_out( VwireModule_io_VwirePorts_0_1_4_out ),
       .io_VwirePorts_0_1_3_in( ArrayRowModule_io_V_wire_out_19 ),
       .io_VwirePorts_0_1_3_en( T19 ),
       .io_VwirePorts_0_1_3_out( VwireModule_io_VwirePorts_0_1_3_out ),
       .io_VwirePorts_0_1_2_in( ArrayRowModule_io_V_wire_out_18 ),
       .io_VwirePorts_0_1_2_en( T18 ),
       .io_VwirePorts_0_1_2_out( VwireModule_io_VwirePorts_0_1_2_out ),
       .io_VwirePorts_0_1_1_in( ArrayRowModule_io_V_wire_out_17 ),
       .io_VwirePorts_0_1_1_en( T17 ),
       .io_VwirePorts_0_1_1_out( VwireModule_io_VwirePorts_0_1_1_out ),
       .io_VwirePorts_0_1_0_in( ArrayRowModule_io_V_wire_out_16 ),
       .io_VwirePorts_0_1_0_en( T16 ),
       .io_VwirePorts_0_1_0_out( VwireModule_io_VwirePorts_0_1_0_out ),
       .io_VwirePorts_0_0_15_in( ArrayRowModule_io_V_wire_out_15 ),
       .io_VwirePorts_0_0_15_en( T15 ),
       .io_VwirePorts_0_0_15_out( VwireModule_io_VwirePorts_0_0_15_out ),
       .io_VwirePorts_0_0_14_in( ArrayRowModule_io_V_wire_out_14 ),
       .io_VwirePorts_0_0_14_en( T14 ),
       .io_VwirePorts_0_0_14_out( VwireModule_io_VwirePorts_0_0_14_out ),
       .io_VwirePorts_0_0_13_in( ArrayRowModule_io_V_wire_out_13 ),
       .io_VwirePorts_0_0_13_en( T13 ),
       .io_VwirePorts_0_0_13_out( VwireModule_io_VwirePorts_0_0_13_out ),
       .io_VwirePorts_0_0_12_in( ArrayRowModule_io_V_wire_out_12 ),
       .io_VwirePorts_0_0_12_en( T12 ),
       .io_VwirePorts_0_0_12_out( VwireModule_io_VwirePorts_0_0_12_out ),
       .io_VwirePorts_0_0_11_in( ArrayRowModule_io_V_wire_out_11 ),
       .io_VwirePorts_0_0_11_en( T11 ),
       .io_VwirePorts_0_0_11_out( VwireModule_io_VwirePorts_0_0_11_out ),
       .io_VwirePorts_0_0_10_in( ArrayRowModule_io_V_wire_out_10 ),
       .io_VwirePorts_0_0_10_en( T10 ),
       .io_VwirePorts_0_0_10_out( VwireModule_io_VwirePorts_0_0_10_out ),
       .io_VwirePorts_0_0_9_in( ArrayRowModule_io_V_wire_out_9 ),
       .io_VwirePorts_0_0_9_en( T9 ),
       .io_VwirePorts_0_0_9_out( VwireModule_io_VwirePorts_0_0_9_out ),
       .io_VwirePorts_0_0_8_in( ArrayRowModule_io_V_wire_out_8 ),
       .io_VwirePorts_0_0_8_en( T8 ),
       .io_VwirePorts_0_0_8_out( VwireModule_io_VwirePorts_0_0_8_out ),
       .io_VwirePorts_0_0_7_in( ArrayRowModule_io_V_wire_out_7 ),
       .io_VwirePorts_0_0_7_en( T7 ),
       .io_VwirePorts_0_0_7_out( VwireModule_io_VwirePorts_0_0_7_out ),
       .io_VwirePorts_0_0_6_in( ArrayRowModule_io_V_wire_out_6 ),
       .io_VwirePorts_0_0_6_en( T6 ),
       .io_VwirePorts_0_0_6_out( VwireModule_io_VwirePorts_0_0_6_out ),
       .io_VwirePorts_0_0_5_in( ArrayRowModule_io_V_wire_out_5 ),
       .io_VwirePorts_0_0_5_en( T5 ),
       .io_VwirePorts_0_0_5_out( VwireModule_io_VwirePorts_0_0_5_out ),
       .io_VwirePorts_0_0_4_in( ArrayRowModule_io_V_wire_out_4 ),
       .io_VwirePorts_0_0_4_en( T4 ),
       .io_VwirePorts_0_0_4_out( VwireModule_io_VwirePorts_0_0_4_out ),
       .io_VwirePorts_0_0_3_in( ArrayRowModule_io_V_wire_out_3 ),
       .io_VwirePorts_0_0_3_en( T3 ),
       .io_VwirePorts_0_0_3_out( VwireModule_io_VwirePorts_0_0_3_out ),
       .io_VwirePorts_0_0_2_in( ArrayRowModule_io_V_wire_out_2 ),
       .io_VwirePorts_0_0_2_en( T2 ),
       .io_VwirePorts_0_0_2_out( VwireModule_io_VwirePorts_0_0_2_out ),
       .io_VwirePorts_0_0_1_in( ArrayRowModule_io_V_wire_out_1 ),
       .io_VwirePorts_0_0_1_en( T1 ),
       .io_VwirePorts_0_0_1_out( VwireModule_io_VwirePorts_0_0_1_out ),
       .io_VwirePorts_0_0_0_in( ArrayRowModule_io_V_wire_out_0 ),
       .io_VwirePorts_0_0_0_en( T0 ),
       .io_VwirePorts_0_0_0_out( VwireModule_io_VwirePorts_0_0_0_out )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign VwireModule.io_VwirePorts_3_22_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_22_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_22_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_22_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_22_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_22_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_22_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_22_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_22_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_22_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_22_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_21_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_21_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_21_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_21_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_21_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_21_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_21_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_21_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_21_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_21_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_21_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_20_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_20_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_20_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_20_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_20_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_20_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_20_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_20_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_20_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_20_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_20_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_19_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_19_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_19_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_19_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_19_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_19_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_19_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_19_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_19_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_19_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_19_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_18_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_18_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_18_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_18_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_18_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_18_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_18_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_18_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_18_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_18_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_18_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_17_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_17_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_17_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_17_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_17_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_17_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_17_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_17_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_17_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_17_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_17_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_16_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_16_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_16_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_16_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_16_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_16_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_16_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_16_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_16_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_16_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_16_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_15_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_15_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_15_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_15_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_15_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_15_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_15_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_15_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_15_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_15_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_15_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_14_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_14_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_14_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_14_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_14_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_14_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_14_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_14_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_14_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_14_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_14_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_13_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_13_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_13_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_13_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_13_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_13_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_13_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_13_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_13_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_13_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_13_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_12_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_12_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_12_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_12_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_12_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_12_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_12_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_12_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_12_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_12_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_12_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_11_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_11_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_11_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_11_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_11_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_11_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_11_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_11_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_11_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_11_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_11_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_10_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_10_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_10_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_10_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_10_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_10_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_10_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_10_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_10_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_10_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_10_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_9_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_9_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_9_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_9_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_9_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_9_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_9_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_9_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_9_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_9_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_9_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_8_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_8_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_8_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_8_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_8_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_8_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_8_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_8_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_8_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_8_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_8_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_7_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_7_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_7_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_7_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_7_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_7_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_7_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_7_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_7_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_7_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_7_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_6_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_6_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_6_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_6_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_6_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_6_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_6_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_6_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_6_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_6_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_6_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_5_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_5_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_5_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_5_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_5_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_5_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_5_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_5_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_5_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_5_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_5_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_4_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_4_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_4_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_4_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_4_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_4_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_4_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_4_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_4_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_4_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_4_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_3_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_3_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_3_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_3_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_3_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_3_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_3_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_3_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_3_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_3_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_3_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_2_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_2_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_2_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_2_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_2_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_2_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_2_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_2_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_2_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_2_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_2_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_1_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_1_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_1_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_1_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_1_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_1_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_1_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_1_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_1_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_1_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_1_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_0_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_0_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_0_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_0_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_0_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_0_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_0_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_0_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_0_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_0_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_3_0_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_22_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_22_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_22_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_22_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_22_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_22_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_22_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_22_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_22_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_22_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_21_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_21_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_21_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_21_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_21_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_21_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_21_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_21_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_21_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_21_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_20_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_20_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_20_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_20_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_20_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_20_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_20_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_20_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_20_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_20_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_19_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_19_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_19_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_19_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_19_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_19_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_19_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_19_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_19_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_19_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_18_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_18_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_18_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_18_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_18_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_18_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_18_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_18_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_18_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_18_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_17_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_17_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_17_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_17_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_17_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_17_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_17_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_17_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_17_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_17_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_16_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_16_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_16_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_16_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_16_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_16_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_16_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_16_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_16_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_16_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_15_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_15_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_15_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_15_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_15_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_15_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_15_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_15_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_15_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_15_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_14_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_14_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_14_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_14_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_14_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_14_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_14_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_14_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_14_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_14_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_13_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_13_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_13_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_13_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_13_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_13_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_13_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_13_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_13_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_13_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_12_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_12_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_12_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_12_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_12_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_12_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_12_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_12_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_12_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_12_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_11_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_11_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_11_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_11_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_11_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_11_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_11_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_11_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_11_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_11_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_10_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_10_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_10_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_10_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_10_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_10_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_10_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_10_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_10_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_10_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_9_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_9_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_9_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_9_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_9_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_9_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_9_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_9_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_9_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_9_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_8_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_8_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_8_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_8_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_8_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_8_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_8_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_8_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_8_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_8_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_7_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_7_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_7_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_7_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_7_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_7_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_7_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_7_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_7_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_7_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_6_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_6_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_6_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_6_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_6_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_6_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_6_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_6_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_6_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_6_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_5_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_5_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_5_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_5_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_5_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_5_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_5_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_5_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_5_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_5_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_4_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_4_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_4_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_4_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_4_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_4_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_4_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_4_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_4_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_4_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_3_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_3_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_3_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_3_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_3_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_3_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_3_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_3_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_3_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_3_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_2_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_2_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_2_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_2_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_2_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_2_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_2_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_2_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_2_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_2_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_1_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_1_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_1_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_1_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_1_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_1_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_1_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_1_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_1_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_1_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_0_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_0_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_0_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_0_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_0_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_0_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_0_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_0_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_0_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_2_0_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_22_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_22_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_22_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_22_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_22_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_22_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_22_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_22_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_22_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_22_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_21_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_21_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_21_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_21_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_21_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_21_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_21_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_21_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_21_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_21_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_20_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_20_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_20_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_20_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_20_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_20_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_20_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_20_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_20_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_20_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_19_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_19_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_19_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_19_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_19_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_19_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_19_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_19_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_19_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_19_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_18_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_18_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_18_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_18_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_18_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_18_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_18_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_18_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_18_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_18_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_17_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_17_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_17_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_17_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_17_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_17_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_17_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_17_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_17_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_17_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_16_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_16_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_16_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_16_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_16_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_16_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_16_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_16_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_16_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_16_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_15_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_15_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_15_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_15_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_15_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_15_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_15_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_15_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_15_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_15_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_14_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_14_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_14_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_14_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_14_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_14_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_14_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_14_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_14_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_14_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_13_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_13_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_13_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_13_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_13_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_13_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_13_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_13_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_13_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_13_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_12_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_12_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_12_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_12_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_12_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_12_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_12_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_12_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_12_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_12_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_11_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_11_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_11_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_11_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_11_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_11_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_11_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_11_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_11_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_11_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_10_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_10_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_10_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_10_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_10_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_10_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_10_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_10_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_10_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_10_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_9_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_9_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_9_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_9_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_9_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_9_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_9_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_9_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_9_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_9_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_8_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_8_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_8_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_8_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_8_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_8_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_8_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_8_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_8_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_8_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_7_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_7_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_7_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_7_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_7_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_7_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_7_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_7_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_7_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_7_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_6_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_6_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_6_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_6_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_6_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_6_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_6_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_6_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_6_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_6_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_5_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_5_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_5_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_5_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_5_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_5_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_5_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_5_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_5_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_5_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_4_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_4_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_4_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_4_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_4_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_4_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_4_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_4_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_4_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_4_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_3_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_3_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_3_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_3_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_3_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_3_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_3_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_3_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_3_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_3_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_2_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_2_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_2_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_2_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_2_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_2_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_2_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_2_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_2_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_2_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_1_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_1_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_1_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_1_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_1_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_1_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_1_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_1_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_1_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_1_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_0_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_0_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_0_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_0_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_0_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_0_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_0_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_0_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_0_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_1_0_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_22_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_22_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_22_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_22_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_22_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_22_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_22_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_22_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_22_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_22_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_22_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_21_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_21_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_21_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_21_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_21_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_21_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_21_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_21_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_21_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_21_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_21_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_20_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_20_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_20_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_20_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_20_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_20_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_20_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_20_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_20_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_20_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_20_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_19_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_19_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_19_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_19_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_19_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_19_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_19_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_19_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_19_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_19_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_19_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_18_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_18_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_18_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_18_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_18_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_18_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_18_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_18_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_18_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_18_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_18_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_17_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_17_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_17_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_17_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_17_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_17_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_17_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_17_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_17_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_17_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_17_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_16_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_16_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_16_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_16_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_16_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_16_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_16_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_16_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_16_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_16_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_16_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_15_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_15_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_15_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_15_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_15_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_15_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_15_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_15_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_15_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_15_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_15_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_14_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_14_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_14_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_14_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_14_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_14_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_14_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_14_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_14_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_14_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_14_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_13_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_13_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_13_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_13_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_13_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_13_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_13_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_13_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_13_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_13_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_13_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_12_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_12_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_12_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_12_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_12_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_12_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_12_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_12_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_12_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_12_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_12_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_11_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_11_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_11_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_11_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_11_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_11_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_11_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_11_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_11_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_11_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_11_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_10_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_10_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_10_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_10_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_10_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_10_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_10_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_10_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_10_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_10_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_10_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_9_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_9_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_9_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_9_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_9_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_9_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_9_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_9_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_9_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_9_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_9_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_8_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_8_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_8_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_8_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_8_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_8_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_8_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_8_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_8_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_8_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_8_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_7_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_7_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_7_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_7_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_7_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_7_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_7_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_7_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_7_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_7_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_7_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_6_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_6_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_6_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_6_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_6_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_6_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_6_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_6_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_6_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_6_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_6_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_5_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_5_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_5_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_5_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_5_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_5_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_5_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_5_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_5_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_5_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_5_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_4_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_4_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_4_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_4_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_4_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_4_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_4_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_4_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_4_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_4_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_4_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_3_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_3_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_3_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_3_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_3_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_3_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_3_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_3_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_3_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_3_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_3_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_2_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_2_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_2_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_2_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_2_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_2_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_2_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_2_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_2_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_2_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_2_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_1_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_1_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_1_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_1_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_1_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_1_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_1_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_1_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_1_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_1_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_1_2_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_0_15_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_0_14_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_0_13_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_0_12_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_0_11_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_0_10_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_0_9_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_0_8_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_0_7_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_0_6_out = {1{$random}};
    assign VwireModule.io_VwirePorts_0_0_2_out = {1{$random}};
// synthesis translate_on
`endif
endmodule

